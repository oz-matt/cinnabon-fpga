-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
eoyIowv5migMojZk2ZdhS1vZUb/duXq+WAPdfARRSmoWsGKx+V5f/vCiG8cfcIKWDyFGtuTqxoKf
LLMYgiL1jgjR9z8mGsj/57dYvzMm9gnDTATvskUqYB1jc4ikL3A8asGngSGjUKh6GJrwmsv1Luh3
3a3i/UGWQZAc2Plx97ml9eP99uTRcC7O2fK3hkD/uvI2cMB1aNCzrLOI/fwt7HeAk1/2zrCBsXx5
3QVFH3vq0tAeWZ9LSUEgDnBz2JLJR0mSOXOOp+V125KOA38b5ArwDS3nqYSZC+6wJTKplG0e8Oc5
A7SpLa4Tc9PlBb8dUPRGsxRVaTxKICfoSGaTmg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3632)
`protect data_block
wiZ6M9dfrYL6J0QmQ+jS//MbDz7jafQeQRVByGNQbw27URk7K44PUJZ0DmOn69fli7bFf8i+KfNe
Ts5jkEdmK0g49L60u/BGYe3Cf4hHF/rfpeXK6cHqxvwmuVgiTzJNuofXzqHiceZKsFNjkRj/9J6/
naoqDj7E3Y0u37hS++O2eYXKOf1gfageT/w8KH0Rr02Z9ipzwuNi7qS8tVoDBk7QjeuzIjyyqzmY
4eozSkStJgPr51b4gRjA9oTPmV7rW0xWDiAiLs+Qwg5jMiVKv0eTwOgsk64BESix54wmmgOalnNj
wXStvOy4WzuEps2dEEnT5QJzThvrzqhYP0Xjm0e1xwAXQoWtl4svfSU5cqUebOMPQcUCITe3rirG
KRaydROPpv3LgaEMQQ035lM+1RlF/x3zq6Auuz5SrRr3MygM9gRRNSRFtUQtFQlAiZ7vNb2Pwz9H
3mx8Ds5ffWFV9JhRjwKuN66+NHrk7xIo/CPkHP1Y5GHXLqyWf3wybGkB4qAFAR3c7nU/lzQM2EEz
0Ba/WQ4ZcnGSBDf4BTDgqcgYgGWgDz5t7lfzEeAld4254NJO2v4ESC+1UEIwNr6ZFQnKk52QeHwR
1HAcTI4eZuijtCb/h/d+2Z/hzh9OLPErDml61rs0G8bQI6yza8wTqdwGj306OuOZCRTpRt4hfR9N
gWM5ncKP7gr1A4xzmZPlm+gedpdH5eXqSkmrPskDG9JAF+r/oPWcX4cYKQJwP+H8Lo12yqhjBpCo
tueGuvbR2TQTUWeZ+/nngajuGTEbOYUWmzBWhp+h3jtFi6PN4UoWPoOg+jeB/gnqR79XiWh+NVfC
SbtgIEYIRbVEX5T3RFbdHM6+VPYMIAbv1MMNe1bq7OEQf0h9QrMDG6Oj+LhawHxpjUDVz6EC5n6y
jB/SOXuCDtgCNiVs1+e1IBMNsZQzb0gxEw8vgyipOE+mJYWVV9N2EZFtxGW8Nx8FjvikcIuhswua
bi6nMpkc0Jlvt097QnOrETHepzJdQcF3xCT+h1IrBl1/RMlmuGCHbp4VXZmkGo1P5XFZMK+VL8dl
mqsSNlF4Q6Rdy8tMqKdtIHE2EZ7Cs3kqMlV6NcvG5bKa4G/8tXC702UcOxsxOst+fMAwxETu4E4T
F6mlz+KKwxAeTn5H51wbN0znKGDihbnPoBu+LteC86HQpBua42BzFjOWrFjKTOaLlvZM+emufmc7
bxSEmku1+HDShSOnzf+CjsgyIX8w5y6iQLsZcxjcixQpNQS5MIbjkyDhRVbZqLSGOFH+LBJqKdGK
9cV3sq5L6iEbA2SUKrZfJVF4Of/T1+SvoG+2Vu7v0O3L/Vn8YyHR5h8dBzbOOqFI0cKNmqm35dIu
MY70i7tCe5Bs7EgnXcEWvI0ic3xZ16nTqQK2bkoJprF1AL4sGzzqT/iXPo6ar9h0MgotDyLLsCgu
U1cO4I8WaUSzqSE2OQMgkdHoJsLGOsi2MrF5R3q639RxUCVFxaFvHEK6KRL43ex+k1NMrGbzFXjk
j9ysG/h+RV87bUplm6gcowO7qGWAthnaqJ/1YZoHBIMTNrPP1LtcQ4EvW0J5mWFeI163TBab4/yd
ahojo7Hq94nXVgSk7r7Ag7lRXNpm3M4KYrJKvQmshUcBsCVb8aHQR/f8+svuSMsB5nKD2Rke1AVD
a9S91O163SzvrZ5lvoG5d3sb3bobNZIhGG1CtSbFZJGMHqO71RnAt4Z/Spa0RclW/dgqsxxjzKF8
3ERFcHDSpv6avNafPAl05BqGQlxTvITZE2DMQa49BoG+cy7uZCd1piPtKf7o8PVZEpcw0L8DcYUw
Ly5D+X/rx9A5LiA2Tk+tC+kHZ17rqBIIXdKZchleV7Cn5Cdykjr7e+FUn5l8IUeLylnPnP4w2OfB
QiMX9cFjuhpzsSxJMUZt6CMJlopc5qIu7MLPjtwCIiw5VULQ52sNtXjteS/mOu+TcknhSfLNnz32
Ak7U+dQL7VwvNddeFoJKZ+Zypccr3247apbaxr+d3KrjfCnVHSxLyuW5iW/0c0Hnj6cHDLiiOea1
mzsZNdHxBEVIHok+j8OO/DN5lS/OqOQ8lz2iTLg+xNysxhigtm4bvgOSnSWkBRadysAsMU13DrV0
u8V35JhWbnkc9r0bCTSrcql/59sp148MhTDJaR+OzYDM3/SiUgibBygJ9zoM3Ht/UaDkguaUj+BT
sReTc2P52AHT8fLvnZUakIhDYcuhtpvtLY/AND2Ds/GioNcxPVAf+f08HsL4FJnypN77vIIUhpbW
lSnVa2bqxnB/D1+G2j55cKfWJoo23eGZ1Igq7cihXgfQwnOLNFoOmuTOwsdgkMlQIZeVwDCF9EVW
+uZkysw2J5pcYi54Wd8KPkC2EljNlafO5viTa3258LnwmEln3TT/4bFaW4h6BTdd8kiA3aK7d0DM
EgSIvh7FJExUsuZVABPexcuRSgxfJfaKfurjwrTlX2evBiKwlgPBnhWMX1qQIc74Poz+6gCk0WQ1
DWoxePtKO2+E4WgJScrVkWMpad78yMgHbBGk/rnhGE6gqigayY5z/z7sHgwZ63/LkGoCn1I2hvXT
JtSF9Lk0MofVmISpOsC8bkWOIDfNjEF6I6f9XOMACxBAuF5MtzwkTRlyxej+G8UqsH3veTCOCSO/
5zIEyjwpoxtIOBvU/nH2AE/lLU9fRLU+2GZEIuMb/SWoOz4/XaIsWP3a7nCxxb6M+36p71l7pa//
dWhvmBMi7BKyN99vv7FfwRdqnPK2o0fuAi0I6iUGoQao/RvEo0fMJn29luNq+7gIrhi4Fzuio2HK
8rxLnEILnhRInj4jcsMWNQtP5CL9xhgFu/9vjRCQyI4FtK+XPwr/Kj9ZYMiVge6ztiuq+0V950Iq
3Fj7Ip6i9y31FJAAIYFFrt83yS3ayepfWCJZ6WKFQGnLhqU+yOIRIbAf9oLnVIuVITUY9cbq+D9U
jAtkxCYhthsh6AN8vNTu9/3Rbrd5kF+JVw8e282oLtswLYYtQJfHcfe5YKj+lQhkvsJMaLtcUTpw
l/6cF0vc3Mwtgaz4IxC6mCJUXYjxhGZSEOC1hps+TVVHv7Y0DmJPy3zsqYXtlPQL7BmZFiWSNEME
uC+B+xR6EoGQKALRwF7h5Q1Zofq+sJnJtuG+dmYhSzt9759oONHm0ofB7D0YGCHV13Vd1MeITgEQ
ovqwDeN8Vnvds+d05cm37mMJFUg75XzzmPdzaYkVM3x2ilHmPkIcCKYCAkaXvrdr8J9g+wkZlKLB
S82Wh8dqk7xBth7Eg0wMD2Jj6ZXKM+8Rdq/7bJd9/fnK1tgeAOdURCTLzyOqvcMUmp41BNnslF3x
BNrACPH98V1ZIve1jaquHCQwQZwNn43/AOVqx87B+1d+mkZN8wVr/E97Kl5ail7vBmxrmFpwyLR7
snZx6gQo6iH+2ljNWa+VrlHp/oKjoTVFVCDYbKAOxIjRjVFz4f6+Ver3ejRt4aGSqEMhbDG8/qpD
wTHz4hXmKr2VHivln2Ho+Tk9ohIlvMUTbo/95+cIh/jIk4ac3G0I0Srkey7fV/wwgm2nUF5b8SbT
jh2Ld+ykOurvHCNzy9BPh90iiG+NYLLr4Xl4OSYLCCgocSXeKng+Yuo4v8Vqd7A9B+pAM1urSuWO
xonrYTXBhCnWmypwqU+aTwfE7bgf/erh1th63cQBYEfeWG9131Buc/R0z2BW5v/3dHpzklZDqxin
Eg0z1FlHKqfjSJtxPzRryTdudmu1qTRxwyN0HcQHVgDHP3N6jm5AYbVfWWf80GHMsgy3qXoq+8rt
d6+lNXcvFOmmAseieK3b5Q32KVWsTJaFX3/n4pBmXkTs5LiKFuquQOynRcIfXnJR/ky4ye7rnsJO
YwwzxcppPwoVpd+SkcSAf2LVLPansAjQQbbNBC4s1+F3K+1+HFezMwtaeZPa4U5bQi8LDokVk5ia
Z6ry4oflntMYAXSPxb36EguUpWLJjDGhVptzHtdZiWi5ZGnnJydOzg1utcrliZOqPprxE3KSlB82
XOLj/LPowRGctWZHg9uFnJPU209abd8uQTSo6YtnAripIDuZZuZM9mis9UPLVBkz55ks/02kde+5
W/8VadFgB2X4Ekk8KUEr4TNOyOosDbkzlZ6JhdzopspSdEI81IlFoiIJQwSL8HL+OBVGd5k+2DfO
wWdSoL4y9DXO9Cz+SLv5Em7oMERnCpxIi5zF/sygW/6oXAQCfm5XMkqFTNXaxCBzPmnH6yEdB3re
oeCiEmgSZF0HowYLlw9EBcLhV1HALtz41bJCAefnyTCSsbVjr8lbKyCkgoMEtSqku84y8K4gRAyl
+aQutzyJMlmRnyCVb6jn7JhE4pLWqyjGem2vxP7JfN8JywM3Uhf0OGNTbkYmhsEkRSOkYgjd2Sk+
d2M9AiD2eoPByzlyJZdoAlMMJ5HTnGR++/y4nnFexD+V9i9yo/MWkwdrOAcl3/PhGo2AvurLt3Dv
YMZQM6utzZpvExHLpYMNfAOUZVi4MAEjNctmJbWX+8iJD3Oqzi8gSbW5Vp1YKtM7gMx52QpwGr4D
R/yzEdV2CD12GE3pb+gFKIShdhWXcrNV6FI8Ci01vMuhZPp8msr/3nUPzzkJnVvuGpidOXAMYUbQ
vudGxddHJ0q2JyhwG2SPYSYjP1dZbpM6ROjOMVaEGunC6Yuq/XBLOfaI2l4ftSNjxIkaH8dR6oc7
X2E28ar7QYZjklZZuOVjZfVAOBZ6KqW4EIIYRV/proSxgZ0M6TSTQQ5hqNs6zfeJx9D7RJZV+OPN
0rZvh3KuabJu68meMjL9YLAcCNXcf/2pbUkm77n/213ccaW9zCbkqY4=
`protect end_protected
