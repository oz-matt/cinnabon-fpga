��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o�q(��O;*�|�%hW<ݛ�!T&��q�T��%�^�|���`�A�vG\� ��,o����?��)��Ba�۩�51޳_��$(��&"�҆��*%U�O.,-�xt��IV~�;���b��c�@�����&����5�؃>��j6}2��I��E�QT���]}u�$R��&�cײ��^�`�f*hrݬ�6�_U��F��9�i�N���Gk,�߬.kQ;��Q��x	�|��X�ਝ����H!p;��l��0X�j�$�o��5��s�������9i��J��+,�M����)����K����3���q,I�Z�ml��z���'���{�V}ʾy;8F�E1���yEg��������o� W9��	�Z޾�@/$P���]kM�?�L��)���%ûs��2*q.x;�-���h�r7낦����?/vj,g����9m��E�w����jpBkA��+��w������y�X���^?"�C7���>���L�)�J����ry������{��wץ�'�>��im���&�A3�����{��aQ�*(��(�n!��o6��ň��U��Q�ʠ���W���Q*��E^�өٮ'�2܍��l2A�	n
8�r�l7d�H[�e_Z4,��W��ؖ� �r ��蒾��{�(��	�Oc����p.�X�c�9S:�&�TtT\ް�V\����>����ֲ֠��-TtC�FdB*Ȣp�Hȗ�6�Ò.��T�K���ʞ ���k=+n���{$V,�꿙B9����Ԉ�����6m��i�t]�3���ZFF}�A���)o�>5���Nvi�Fk'�b�lL�=��@�c2h�-����Œ�Z�Z6L�]ی�Y��q���#����)��u�-&�F)�fij�6ʕ���t����)2��o ���<�d��B^h�?�x�7�[=���p�HP�Rm?1t���.q��F[޺�2�F�����e툰�A�I�'�ϹӳHh7�tI�Ԝ�Z���O{6dw�=s�[�` 1��]K|�P)og�P[2=N�|0��
n@V�Tv��"�}6#Wq�	�����6ݣ7g��)��T������l�gM��y�`D�T�
(`�i�2�"G��!�/��!}�=��e�}>��'�'j[=;�R�6��'uyÕ뛬�k����8�:�*�+!�<��p��_�z��l�y0{A��s�U��o��Y�����$آi7$�/�
(T��hjr��Ԁ�b���ob��cHO��������5n�)���N��dy�Pr�#���n��3�-l��tJ��*�T)
0��5I]*'����~�	0c��B
Ȃ��<[0i�Mk�OwD5��V�ub��\;���O9�QR/[!{�T�I�����Q�o`Ū�0Pn�M0�0Y���U�ITp�n:���vHǄ�L��=�rK�t�"{'�m�<�?Gk�C+0J^�V��Y'SR)�Lβ{����MǇ߭��37�e��櫆�C'�|sy΄����g��{ܜ��!Q��U����N�H�?�j���7]!�.l�^�qlg�lu)�@����P��_���ֆӴ��C��RVQ�X��>G9�t�+I�7��DCe�[�2G.�]"�
?�;�C�z�d�S�3�e��g���X�G(�������ƅ�a�A��-j�1��c�e4��蚌�c�szA	C/C��C��6�M7�/(i�Vx��X�d� P�i��uI���?�m�|8�X�[LQS�W�&+�"1��v�������'�܎ߢ��Ƴ��{йS<L� ����=�1�`w��U��~���kᤋC�w�'�+�X=�u`�x��=9I힯��/4��N?���&  N��6����KȥF0!Mʋ#��7(gJ�J�8��� �5l�7�:�(������ӕ!6fL�(�Fz��g<%����X}-3�ޏ�ۓ4S�^��Ƴ�J݈����3�~�t�m?���n,H{���ts{��`<6E��҆�	6��K^�\�żt�A�?�D���]�y�e��\��qzM��yWH�JmЏ3��,w5���3�F�P�$�����X� {�d���k^�̝(.29��]��K��#�
N�:�ēOxu��k����,�is�b/�n?N]ǃ"�ݦp���__	յ�H����L�9&����/���P�i��ԩ�:���%K���_�tU�@��uo�`0�!�r:ӣ����(��տ�H�ZH�B�S���ߜƩ����OR�X&���j;PuE���{� �� H��0�q�����f��
BC��0WhU�F��g����3?�<����;s�c�s��kcH��G~Eu�����9���"X�+��q�k* ��Ǆ�/�d��f?� ����;�-���{1��L�֖�*h��������~�Z�m)u�Hѷ��[�Ф�i[�S���k� d7��u@�����gpA����[�x�nI^�Z�~�ڝ�1��{@�N*�ޑM�1�i
�N��E���a5Ǥ���-�^U��C�=�On�Ī�_ȯ�(o[�=��W�����T��'�t�C�CU�xT�~q�o�i�?FwS�d�Bf1_y�N<���%i�N�7�A,+i"��	���]�Jƫ�$ao��hg�t�O_�e"�~�D�C1�TûK?���$�+�1�5�z�"�/�#�=ͮY�&'>[d����	���4��W ����4�+�<\މ���h���%徥��_�b��L�CbFqxr6P��G\�Mg )W^/3�a���ӈ/��vU6B��%-�y`���9�n[t����f#�Vh@5����uEW˄^!,���B����g;"�yi�n�-i����=�h/#V1�z9f|dq���`d��[-������S�O��R��̉a��R�6���� S��ѣ�����m7e0�%S�3�ݘ�:��׽s]� �l���(㶯
�_U�{`���A���Z-s�w���2Yemb�"��"�j2C����.,�� ��8� �Jƽ�?�#�-!R�`��|�F�ӉyeHK���Y�Μ�'U㱞�N��2��)���85vJS&f\\���A�GwWŬ��V0�\1�M��HHY�`fl[�P6��c�G*�8�\�)2��J}EXa�&Ix�6a�]��0�ո�/��d��>���\c�j�����'ұځ���r�b�4gv,��z��X��ws�z oD�V�6mx�aIF��=n��x���?I�rEY� ��Rf-vd93x�����5����8)�Y�OS���S菦���"�?C=���eh���)d"W�?�-P�i�q���xr�gɧ��s%�12�g>�>r?o;6u{���*6��� g��y,�;�b�J��Q����^b��Т<*N�|�Ť�l���,$'~�(v ϱsR[Ť���锚���,��"��Aj΂�]�9�R+B�Cx|�wLlN��]�k�$��	9�Οt�!Q4]���LFC�(���\mf
�D��7���`|>����S��2WfW��DA�3��mh�d�ޕǂ|*���b��KJ����n�a�3p:ձw>��z8�TO�K2�K��Y�ݺd{�`��[ω�T�����C�g��hҒvJ��~i�j�����ԅ���|��/-����	���k1��V:�΢7=?� ��t��R�t@'�zY��D�U:�#&os��l��r�.�k% -���P��.����t�4{��4	�C0���u���X  *,Í�t�=�ӧ����.<eqdC�=,�|I�P.�$�%��Gu̫�\�	�E��\Z[�Qb�|����|�.V���~Fϑ���c�������3q!m���KC��H��w���e}n=<����7���k��m��X����Y�;�)�����B��1���1�F��믨�<��VY�������S[�o5?�A\��L���1��V�#�ӢEp�n�q��FQ|��/4!-���[]�k  o�K+z���Ť+��q��x�%Vl��*��OQ��6��׽ D1r�~ӗ�)U�,��W���5�-ݏh�f����/K*�_��A�ZÐ����l� �����1i�Q�/^���q�Nα��S�ȼ��#O2�5}�[p�LT���!��e�$܀����y{K�}4	�` ty������g%���P�	�}AJ�	��WWRS4.U6�&��G��yX�q��:Ds�7�f8x~0>���FҕP�lX�p��d!�bh�P��k�S�@�Hq�Sv����TRT%M��Pa��1m7纴Y�xSX�m{�e���r����G���C�B?�ɚ_�C�Zx����l@b���!�
�#�]}�X��4����o��.'�XѨ���A[:F�/��Ӈ��ݵI�X`�����9���d:�3���i����,��E���(�,2:�m��#���9��o�����R����@�ŷ|4�=�yO��-�f���6�C:7"U�8Z��h��N���4)Yc�8����I4�l����wD��Ö[�I ���d!m�����g>gy��"�PMv��t�"���t�T��$]/)�m��G�����K�C����J�h6/
4�QA<�F�[+��
�����I{w
Ļ��4޻T�>����̮����u���cπ�B[_��*2�y�+`b\+˘#d �O��S`5k"�gt^��?����_C�o�̄�:e���	�"��^�m���;��Iς��	�=�1?�Cu8�a%IxA<��Yo!��A�F��!�b�(D0$F���Mn5
+PM���0�0|����V@�T~��$���{���*�OMN�D�e2��tpo>
��?OK��B"�l*��`�{m�����,��6��:�g���u�K�!��d�6������� �ʯ��}4��!-��%���N$���*���1�0Ǜ�9��U��,�P5�v�c?OH��ÀB7g�N����bC;t��%>6��_����s�(V�/!9	��)6]��M�`o�?=Y_i:��);	�G�2����H�(eE+ՀS�����*H��c1Ql�e�ߡ>YP�Մ���R�LUh�M���E�`�S~��a8b-�[��ߔ�$�6�m"E�$U�T#�E�h�1�'g�AV>�����Z`g�vҵ��v)/N�@&^y%��rQ���*�Ʉ �^*Ė+CH)�G��ƹ���k/�l�Y�$�6��ϝueO��p�b�q�!	V�v���	jʾ#��6%��)��∏��Zx`�[�oU�oL�4���4
S]�d�q�H�����H"�%����5�3=����oga�K�W�u�5��7�;'����[���ǝ�|0��ub!|�����4O-X<R�nUF2w�>�*i�2(q�}*H����Qڌ؏s�B��L��
�qZ�wh�����屷��so��5ch�/h�d&��@2��l"�y.���tᴂ ���L��wH�����?�M{����:7U���s���5v_�$�����b�g�/.J�~12�x�*�{y�g6���Ȗb�U��&�rW��fwJ= $�R��ܛ/"^����4�4���ce��Wk�aP��R�<�q�lQY[� #���?���U�u�,�t�d;;|�ذ�p�f����M��s�՞C�H_6�O����MzT|yf-_Q�K�.g���K�pP�t���N�:������bV��X�l �w��������;:�G�F<�I"�g���<��tRv�*�k3���?P���;*���s���2#��29}A@�ت���M����\��/��0f�;$�-�q�(	5��KR]��]�˝���cK�����NP��h�HZ!���@^3��K�/�ͥ�h.	�U�i�K����Eä�������;Z�g�Iwj�q�
�tJ'�A�UB;��
5���9\(��|B���b�9��|��#AI�=���D)[�͍�y����?��p��s$ D(^y ���\*M�	�6Çv1�z�멆���ނV�$�Շ���4%����M	�,�,��S��)95���wA�WW%�m:؞O��G�۠H%�NJ��ػ4�OQ{X1,0��B绝0q�n֎sA�	u˼��>-��3�;��e1,Cr&���9�G/����k>�ⴛ�Sa��6��+��D^�����r$�y�l��u�q��3�:iTƓA��/��݂VX������\"�.o�x�$��B��e�!����Qcz;'^�,��:�M�n����E_
E��ƫꈓ�6x^&���I��W(�ǹ�2����W�(�����8vD}-��~��Z>ᙑ̞{���z� +S4xv�9�2��U/#]��8�>O�h��%w����B�Z��	>�Ͼ��S��1g�oF�/EI�������]=#�^'g�]�U!@ Zd�]W���8 �lP,�1|�:�\r'�y1�� G%0چ��+ρ�AB1@���� ��V���ܻWaz�l@%�et�Ys���d��<DۥҴF���c��fګ�����}+n���i�X��W9��}��n]��	l�g�^~���}f+.q5��?��X;k_���O���j6hab�h���r5p(+����4�F��Z<{�ua��H笪����2����Ն(u�iz1�nDLA�O�R��b �t�*:g^���3��By��l%;�&^�}G6ID]��x �d�	p4�	~��;�l���A��Y��c��v3wC�lυ��hG�[�&I�`G -AGՊ��
�,�s���<�<�g�5�+�7���6�� |WMFO���EX;�%��g��~��'�:d�52�HE��� �|p�1�1�u��9:��	6˭�S)�_N��N$Njp�:�]�[-���P���������(?�Sڷ�NhZ����?��M�S������?;�(5�keX�ƿp~I�Ϥ�/�Bu���N��w����h+��J�,)�sQn�ژ᛻�^:����9��sI�(GY��D��2 ����6�FwQzu��� l2uZ�����Y�ݙ���x�f;ϒx�״����7:O�G��-A�4�Zkn7�h����}E�ĥ�E����)B�Ur��ۘJ��3����Ț3�П�T�H��K����������R��̴�Y�޸���kg����\�"�n�������;A�HY�`�\B��6-6�zEv��)�Z�j��ve��Ļ�&��{;�6��>,�����~ Ÿ6�K�%6�����x1<�6�ڐ ��­�]��Y��P��z*7N��v2��D~3%0�ݴ�J�.z��\�W�O��%ry�����'\s_r�mClU쿦�$�!.8���V�8X�>���l�p�א���#�>��H��6$��"�=�W�k�����0U�21�C�{p
�e{���B�b��įsjǯO������E�cue����4D�V)�;J��թ@j>�q��ΐ�2�N��t3;M8�/��P�^D���Bvz��B�W����"`(�&���ʭ75>����n��k������4�ı�N<�߬-��2$�tj}B}Դ.�HYw�q�.
D�K�)�TW��҈�)���$� ����r��˷O��_��/���������jS+	�Fe�S�����t�H��- }e���٧���Z�zC�
�o
�\n	����N��Ԡ�^��cp�C1R �,u\�����T������,�Z]rT��j���G��̢՟�%�f�ϸض|Kջ!��P����[�;�7�*���ן�:���&����-5�Dr�M ������B�)[�rt��7!��
�-�\����H�'e~H�hױ�>��;��+��P\��7��%,�<&"c��"nHy&����)s4�����gI�D�rڍ�8.4��PW����`\A5\'a_��,a̟_WF�r4��ǹ�z�k�Չ��~K6�N��Wco|�V��r����Ps���@a�����ji��ENDk3�^I�-q���i�H���Z'�/�;S���b2���d<V����jA�$����;�T�!8�X�x���� ���%�J�n��|��!*��������لP��|!b�� �<DQ�rM4y��@���W���_|�P��󙥅�LS)l�q�O�G�`m�NIi�t('2��hR}`�t��1�餫��W�����#(OgZ���`�tZ�J���~BDx���&�?��D"d�,�->������1�(CE���ki����4:�P)O=�`�G�B�C���Nݛ�X�V��i�:=�{����ge-R.��İ^(�YԗnXZ�v���'�����<z��j��D��Q�/��'M�~���Kց2L.�L��6t���d��M�]��}�7�Ҍ��86#�9��O�p�C�7F������)�(F&h}�xd�P�\�(m�ukZj0�RN�G#�!W���	��{Rt�c
�Z�1@��������|����[���� �f1�	g���`�p��%�l��f���T���~T��R��>��;��w���kІ�8�����oO(7��!� ������ ��=��xF��!La+D�����xH�糫u��}3o��f��1m�#��U}�'���9���x]jJ���,t��Ȁ=Ye0�	�-�cRd���������[�����UcyT>9�z{����vDG���Ra9U��U�e|���u����Dߚ�ㅫ���!RZ���ț�E��40|;�]�G�/װ{���G�a|%6�m켨bѐ�|�<�����Dw�A���p�.��@���3�N�� ���H��z>3�����s/
?�����f&z���y�ۦ�p�M�4���:Y�ͧ`�F!�:��S��j`�d�\m�9]�v��;�������	��E\$�Grfu�x�=T7P>�wT3���IЬ�jr\���]�>�y"�T��d�Q�cɕ�ܒS�Z�Ȗ'(cL�����c��~���@��۟ǝ�S+�*��I��6}��h�@���_���m^1V��� �>/U�,��:���9r�K��N��
2�>|e'3���O��S<!we%C2!V�8Z�nŭ!�n��3���x��"wL���ω��R'1c�����2����t~*>����S��;��L��;�9H����ϛ�3�R�vO[��h�����v�E�չ�u�u�O�Ơ�f�J�1��A���&��}_7��K�'W�:UBǠ-шs�O`�!��u8��� �W�����I��F��ʴ���f�.���;�F�p�����>��j7��?���$D��8ݼ����W��k��AM<�� 8���<�uX"a�s�����3 k�#Ϲ!
;/w>4�t��%��^e!df�C��Ot�CwS��[8�u׿)�n������z�K�MLR�=+t��ꯋ�%��B��IK�Ȁ9U�Z��)t{?�:u� CV�{��.cV���N*��-R���Q>;.J~�{w��O����tfe�T�+�=<�F'�C�y�Ϻ=")��O89C\�*��R�(���1����l��T������m!�1 G��.6BhDy����$l�;#$mJ��{���:��cK=��CoD�J�~,&%�"g|UΦ���y��L���)B����2�/����:�yn�)Ŷo����r;=����>�ܒ\k��!�*(
y�k%2QM-�����;�S��:U	�nɺ�չk����QL����F�A<�o�g���n<KP�}|����5@���X?�p�*AoAN*�'�,ޒv��w��pМ�<��f����U�צ<��.��gV�L��Db��8N����V"˻d����W'?ў�q�1�Tg]�)�HG�Jf;Z����YN6lu�C�U6��I
{�G����(sa8Q�=���������I�Q�ue	(��ƈt�RCn���}w;
�"oϫ��>|��8m�J/�O�Yl��}w�;
A ��9N�U��e:��Ϥ���d��FVđ&�	;}�31��N�h��!�\a�TP� C�eu�^��9�ط��ϩ��xl�Y�^9�q;�A&I��~L��0��v�'+�zy��o��x�힞^�����v>n��Dg���ӭ5��-SX�̶9���d�S�!xE�+1����O��E.�կ�
��G��(� b*��	L�5���e!Y
y�?�����r�BH�d+_1#9\���B�ܙh���ۯ���#&�L�0�u\���͖���q���a�ҡXY�1������]��˓�i-���5_��V�\������|�H穰<vm�:���0�p�Q-�٢�}M���\�4Azj���}��QH.�\�տ9�4��FF��e1S�*/���>MF�8�4Y%��{/3�������2�V�Q�Xm̦�LH�{B�iK��%:��	�Z��Vd��gT���*���Gg
!gZ���rn��ۍ����q��w�W#�y���
A?�"E����kl5�#w�W6��� ��uR�6S��$�����oJ�u#n��>>���s{4���U�.������җ�"֣zRav�m���N*����u�z����>VƐ<^3�s(��D�J��Г̾�&6�ޢo�qBL^�#����Uϯ�oS���ZR���n)P�:���`r��0OL>Z�o²&X� ����i_�R{[���_�F����(��3�vt׏"ұ=;I�Ԏ{��A ����~�OUa<?/�~>Z�2
�p4*^��#&#@61`D<{����iڕ?�A��P�tG!Z�^nU�G�����I��*!3�h���F��J�5�(��n�Y�ge����+P��/��{��l{����-��x|��<V��zT{�ZQ��(D5s֕m�*]���X5�Z�c*��Cծ���+6ۀh�.�Gl�Y�Z	�{�u��?��w I)��D�*��r)]���0�c��L�P\��Cwk�N>ЃQG�>�
آ�,H�Q�ر�� k����Ě��(���i��)�}��dP(,\'�SG�a8�6�>��c��haTҠ�'�偉�I{�j{�7'"����r��'�?:\���/���+Ό��R~�p&1�h��쇩�CW�೑a�I�iFQ����=?r�ؙl��x��_��ޥDV�)xT�᭄�C�LR��bZX'�B9�Bɮ�!�T�FS,�Uܢb:�� _6+����b�q�U*J�)>�	O|",Ђ�M�����!�E��Þ��������K��&�--d\���� b�d�����#����4�[	�����qMIp�t��2����w�UݘOj`�D}n��2��"n�@�2'��u�8�D�݁.s�+��Ѱ¾����ĩ��B"p)Qh� E���Vč��2!� �����S�5,�DSt1!W��߀��MKֲ�~8z���6�\0+$mcl��7�ö�D8+)Al����y0΋�S\�A�N��/�?-���nz�˰ͫ�MzzE-�V�r�������\bk���=##�P�� �.�8t���GG������AQUM�T��{�Su:�eo���V���ﷹ�8LW/Ϊ'�Ȯ�q�MҎ��
� TJ��B�#wʅ���sZ)����S��'����3l�u��ě��aHQ�a�5���Ԓ�h9�Єo!�M�D+C��tBm+�(6U�����|*F)��Y^�c�$������f��Q$���
9 �������.���O�7P�$�W̧ת�:�e3\�y�5�Z�e�'z���m>�����_���FE��0�{_��|B
��jy��E�D���w.��f��S�sM����`v�6�pǐ>J��E&1p
&G��q:(�X�aZ�^������nL2`P@�-=���)8��d�{Ee�o��`K�+�h���8�ʷ��D
@����T�k)��9@����`s��,K���Tȍ�%����b��ɧB���d`�����J4�8[�[��T��ḑ�?
��Ou��\P��$�!_��hͼM�n|a���c1w�z �̷�2��'���r�����s���o��/ u���_P$����<�	Թ!3P�����(sqw����@z�@��wo�_�JeI��4Zq�+�S~�>�N����F�'��Er�m� \Yk����Z���+mjU�/� -�ul��I�a��X���5�*�'d������[Np��h��@��^@�,�~�)D��8��r0�7�VsM��:;$p
�"�	<�ڂ�#c�=�Sý/� h��_N6Ci�=�Cr��g��I�<l�7�r&�_��l<i�x{54�3h�������UpB$ˉ���)����eP3���ݢ;�9x,���3 ^�"��q�53)�jBO
H��}��0 /OJ��T�^Ȱ7n�^Ÿ[���iu6�������d)��қK=��	G�L.=5�-�c�����=�/���a�w�V6X��y�~@60�/�･�(��Ŧ�7��&I� 6V�`����`#.x�C7iQU)�v,QOi�z��PCF=�O�{#PWB�_/}b�
�-�����{.V=&�_�<�p;w�R0�WO/!$+�[>�R���h���g��*Ko��;@����ؒ4Sג	M�Lb>�B$��Z��������L�R���������o����tޥi6��8]�T/��${έ�a���E�3���t&!d�.LM��zp�%݅�������ƶ�W�}{��%A,y��B��u�<1��w�<��oa�!ԫ�������ö��{*^�AQ��|���gO+�����%6���?�Ȑ�X�L��&���zd��X�<�|�\�<
�B��O�	o6P�UĪD�p�P��d�����t�F��T���Z�ؙs�&jV}B��	��m�c����B���>�J����P1���q�/�Y�������Z�W+H����ĭ���=��|����O$AwuJ����U��JS��Y��bމ�]�\��Z���O��T���0V�S����3��-G��l�3.a.�w�0	l�v0�-BM��q�yDؿK��QS�Ƭ��w�}�+]Mc�s�����	jw��;�[l�&�ׄ��9]��>i��d<�d��9/�6~T�`%p���V���>W��4�8��Ost���ƈ�{R
��g>�	��hY�M�Y��Sc����{���NǶ�{�
���G3�Sj���/P3����2���g�a�H8	'����Hk�?t���M�iT�^t�2M�3s�7N2W�u��#�����?�=5��%����l��y�mÆ^O�����O�v�5*���_�fs5���oށ&>��7�ɮ�Eèޚ��)�e���iYՕpJ�'�hJaX�l�6�@)g헞��d\:l���)v�
�T��u��L��{/���!�_�q�>9 G-�_����0�s�[�d���*_p�7
b���&��ص��d��:��_2���EVM�%fzC��� ��r��c\ݦ�8�)�F <������芋r�ш��'����UU��y��6oրU���9�4��Mgn^� 7��f�*���ƾ���������*���u�\�����L�W�c!��^���H��ҪAeK�ڒ��k��KY�Ϸ�^�4\x�0VYb(H#A�����1���GNm��7J�3	2���O�a��b� H�#L�I�cFr,��D� �x��y9���j+��9��ծ ��j�wWC����
iQ���S�a�d("���=����g�0\`��jӠg��D�dvGus$�SO�p��`��]�\���E�:\�g
��
�]Z�X�49}���9&�Wρ�	�ʀ�m�<�m%"�چ֍�64���>�m��ɤ)XoCBTG�ɀF�[�o����qM��1Ԛ��$�2M�7�^�f�� �I�O1>tW˾�Di=�a�<ެ��)%�"�=P���R�)2�G=���)-ȅx��Gc{�/ya�]_:�#S���.8��Ou��0�0b��@lU��l���<i+���m���O��1.y��dBZԜ&c�@�a�]�/��V%��y=pv*��G�o��WE_5Q��ܱ�y�&�m����`"�<��A
jӎ��h\>\%�;ߵ@�Y,<D�.���Ȟ��ѽ-��4�b���pG��|K/�3la�^���_F�@(��k����~�7Ď�~�b��/����Y��'ܜ�4�@.�L��%�CT�v�`u-[�W1s'��Oc��D[
M@�?ըU�q���n[�Df�m�u�s1N1�nE�Uk�pU���67�.c�|U����a��x</�2�M�*���0�sI�s'��֐X�j��Bf�o��"�/c���}eEE7�/-��L�w-�:��]N�?�+�Xٳ�C���V�
�w������Dc��.jBh�UJzƸ<?�C$QZ�Q������C�eQ���P
���m�cn��!���+>%���4�pu�~ow?���L��Z�<���/p?H��9�W%����B�Lmx��úi`FG(@�mc�'$�{�>ӖE��&ώ<=ja����f6�+�+p^[�l�O�3��Z�ˆ�Y���rO��������0SpHX6?��x���/��zâ���s`6�V_D����`D���z�w�z-��h"��t�Q���Ғ������@�z\��tIMB���Rxhi�%E�l�
s�F��[�\)�m+φи��$�Φ�:��s�g���@��?u»�*��KRALl�c��iA���d�$��%�@�N�ɔXē��׽���y4K'gb#H�4؉���箞��<��"�1Ύ����'��
�������G<����Z�
��s1]���x�j����ؕ�o+�UW�" �b�Q6ov������[����:Κ�Vl�0?z,/v �p^��"b�D�!+ɧIėh|��4�KZ�d�'�g��/&��b�,�6���� "���D���P�ٵ�Z�1��x!9-S0�*5:�"_��@Y�s0��2L_�5���O�Eo^>�"���\�{�����6�m�����<u*�3���,m�;��B�Z���JM=�������:�ء�mmn����B�(��C���,���r��u��]S1�.�vlN	W�k]��Y��K�(�/p
�w{�5�+�Fɔ���$e�t�z'��?5�X��1����,�o,{��bc:z��j2&^��1n��U@}m9�I����@6��}u��g����~��?�1;e�%�5�������5��2G�[�!6���Ht��J�iƜmM��<G��g��.W�x�'t�vLn�����3�ʍ��
P�.�/�<F<G�l.7�%�3 ^ERo� ��dg�ʒF���8|A�q�F��X�^��T�aO�{R�'�z�1G��b�R�1`=��h\�[�$(_�9ggBF��~��>�=k���{]�%pLM0�$��q�zt���9I��T�rY�y4�� O�%M�L��͡&����D����w��WN�H�}�����ۨ�:Pk�XNǣ�F����TB����=��uc�w�$��q
Z����&`�^�ke�@�����Q����ڐ�x���s*�` h��-�ee�gȚ�h�$] �GJ�.���y�=ze���"�B�M�=�.8��q͇j��SQl���l����Y(N<0���l��˪�Wb36�wD������A�7B2S�N�������߯��h�L���	(�}�ږ�tb 3�P��WT|l�"��!&Xr?jK�N����M��T�ѮL�pzD��d�����a
��˿)� ��;�r�a֜�[�|�s��16RC0����*h��҃����>���^[�X(��G-�9�}7C]��Ɏg0�E�"Z<�x)&��Bv�{�U�kuz����c�\~�8�YCJ����K��F����wu��9 ��faG~�K0 _'<���1E����ቆl�MΜ���Ag�f�YE;�m�����A�xE��L�k����uZ�8 �#���S���[m���Y��8�+����yK"�vq/u�w����[@h<g��&Բ��ҷs��G	�[逾��IE�;t��֔����t�L���E.A�%��cH�X����� [O�����@�Ɓ�F��k�t��x��\qm���Q>QX�T�1F�\߆6+�U�' Dy�����+\H��{��A�NOo�`Tf��F=zb礵�+AQ3E���왥�ĐhA,㺎�h1�dUf��:����B�5�H��4�z�����<V"��o�Nm���I��̙���	J�;Q�����o7&E_A86��R b�ݡ�+8Kih�JmJ�@[����JJrn����+�pW"!��^<�xL'�7�l��t���0�UN���2\����݀"��G^�ԝ�y�C��h�o!;	N�L/yGSƛ�=rb�	��nۘ���.�&�'��?Ld� �;O)���? ���!Ç�8���xB��X�B0°�����4%�-^\��a�/��L4L-a�+V�^�jg~�D8�; ��1�8۱�P�3r���� ��/ڎ��ʭ��G⥐���>0d�`-�&^�� �|F�T�ԭ�[=����T�ފ[���zs�1�B�&-���N�C�.���MH�o8pp�ܧ�Q��K�4��'�+��փpt�g��6�S��UΕsM��`���Z��U"ƣ<�q/�8B�5�+uHuo�6�J^}Y�±A�3c�C�R�Iuxn0,h;=�h>����"å�0fp����&.�	�������އ��䒭��o� �H��!L�)���#"�(�\"1HMvLƳ�k��ި���%5J<�bdU����&�E���:��)�9~����*�2���iA�;�ce�����_&�7@�������HTa����vV�>�跃=g��U�b)#�.�����u��Y[�<9�v��1-����qwk+��zn�~��xXݎp�"����!�_��GS�<Q�;z`fZ���w��!�O�5<�dU�6�'�"%W�鹉7I1��fƵ���}��Ts�+N(!�b�<d�yc��7�F�d��_��(��n�̀���p��/֋�]���Ԧ��KL�q)��~7����L��w*&J�b�铑�s%�52���O�����v���?�v��;h��̾���Q��ή��7K�1��T&�ܺ ) �!Q�/�yS�Å�Ah1��/���$.���z}�Qm '�j�ғ-�뎮�	5M)�x;�k5���&�x+�*^�=��o���W5��ٌ�;>��Ǻ�w��� ������C������)�R�:�<x�P{���^�d�%��h,�]���%m���nr�a��F^2n�v��{LK��]&.AJ�ӈ��<��+0.��o/#��3�2˦�/�]`�5 �S�I�H`��Tk����y�E�=�M��]�1L-u�t]���qS�VN�U�+������	�*��2�+J�F���3u�#�#ĝU^�չ�#5{�3M��p�&��	���"x�����~���k�S���W����I�F@W��z�X����b�e�V��2J��.5q��T�|���9o�a|��F�����_\*(-'j2Ǖ�{���W8�qӺȺ�"� <��}�_�5�4��?�|kr�	sK,e�}���q2^�돮�8B��8 '�‶��D�W�-�r�0ٛV0�zc�{��îaATxq�F�L�C�$P����vڽ�,sP$�U�wcG2{��_>�+]3vnO�G]g���+��؆9Dl��@Q�'Y�w���W@?�u�U��Dwy�����9PԘ�R��Z�Ky��i���8u�X,r��ȮE�ӊ���w��:�=�=\����Y��)?��Z�wʋx{�-R`;���:��������v0ñ��*؛�<��nq�O���I�cg��rCr�iNժX.V�<��C����dp���8��\2c��c*>ͿU^�pk>=L9Y��=�)Pƛ���C ���EP�-x\[�ڲ]�i�v��#xbBez�\�=#�'N�У$� ge���P^(%�Go�#)��Y���M��E��<]/6X����������`�s@��A�@#�9WdOF�`w!��3~����ʜ���x�i��|$��&o��A��>��#� [�
��Zz����,��i
�m��_0����_�ܛ0��_��n��3z�̳H�� �z�o
�it���R�ՅVh�����O�*����n�訽W�l7�yp��rA:\'�
*y��3(�{|���Qoh���ɲ��D	 zg�����ۢϘ=n��y4���$�qqJbA�J�|��0ڱ�蘷�Q��ʝ���t!���� �������(�_�F��*k Z+��U��4�T�4N,��d�!l=������8+;r~�v`��|"���|��U�T*��w��b��h���R���|���D\�ٕdQ ��"�����h^��Ԍ��o�
�\�R��~����1���ц\�@Y�B��#����wG����CPR��T2��c$b��0k'fq.�F�H�_�|�|�F�%��Z?>���+7/�;��\g�����│IL��v�x�:r�0U0 �!%Fy��k�`~Af���_-N�t��0"o�o-��w�^łH��x�|і�~e�Pwu^�c���a3��kG�T��bƸ�}�­��L�:>�Hl8�`�t�1,Fx�Bģ\��S�ͯ�RAѽP��	��J	�eƍ�|�].�E�Q=�<�s_����& O䔁�������Q��T1hpH�`���>N��]�4�,o����E��C�_4^��c��3]ݹ[�FB)���3�*^ߑLB0
]�h�,�����W�f}�9|�t`�÷��@Ju&���?�1�봂Ո��Լ�����P'I_���Nӭ춃K�'p��1��q�w��c1,��Ƃ��f���� ��)'������ˡs��ؐTU�%s�X\ !k��4��Q��ȇ�S��<���$ 8X�m0��jS��s��c���(搴'��Р��u�7�W�W�fv;i(C�����`ߞ��p�6�C�~+�8�]���!w��͘����҅�]ɼ �b1c�� v�qKpNs�I 1��ѣR,�O�R��r�Ka�	Z���bW!�U�=�fs��dRWL- 쀪�+�vwȤ��!.�
D=4!��۠�:ڬA
.#>��C�=<������їVX$粸+|!0E�r0 �O�3�Qڋ���{�޾�[_���8�-*�[�G�Q�K2�h��>Z]q�jo\���n�HY(�s�|f�hw���L��Ő�	�^�y��r����_�-�F���!��Kͽ�!4��Y��K��z��w�hV��/�U�J��A��P/�:��"��꿓�(H)X�n��FwT����9'�Ȱ��	`3�����o5�@��h�����\���B���$%]��]"T�_����`�Z8Q� �?�I7c�so�ݖ��c3�@�k��@/ �
$��8����9:�Qn�FI?��bYE�d![���ӓNp��K�S�uÖ�mg�9��Dt����Zp��o
�u��ԟ�;��K'��E}*��}X�q�w�`G�u�[������)����T<G��m�'xbb��Z�(�&��x���b��;�_)[0�<���P���ژ䗑@��xk|Y��q��&3�x:
9{f<�&ѡ���		������7�:�\�^��A0Nm(մ��n�Yݎ_�+++��V9,�3�����%c0��dPz;u�}[�TY�4�/Fu��@��-�e^��؈~d?]n3]	;˕6�f1l�8�#�ymn+�Cd�򎥖ߗ��&Y��|j9X�+-����{C;f��tZ%�e���"<k���Ђ��F�]�q��B����iqs߸h���!���s����X�P����fؒ�<3��Q	��d�г�����z�����E9�]�$�k�'�m����w����� ��F��DtAR��Qv�z}Ec��=<�>Ԯ@�����ns(|��DcQ'G������h^A��p���~�hwDBƆ��(�7�˪$>f�bQSĮe`�8������7�.�z�%�����Qz�홄	G�H��X����$����r��s�gTt�v���J['��օ
�;�dO%?K�����K*HM1ڒy���S�f*�i�_���w�<�|�ǯ��U�*D@M����/*ħ���'L�k,�Bx�=Y���hzY��Lb�wB��A���e3��?feGnE*�JA�T�p`�#�	;���㼈�����Xn��=
zV'���������6�Y3��왵�H?@��Y4i%��p@���~�����`��)�������ǜ�H.��=�����r����qEl~���C��T�Ox�L9��K
������X�GL<�޳�Nmn�h�l�(�"���T�����U�T����8=.�(s�oBJ聛�n�QRC�T���Fj�X���=H�c����O���'�.��h}|��'d4���u�հ��Y�Z��G3ES�?5%<8�ƳTs��>.�2>0���׾��=��\7*8����lh����
<��)���s�bu�FW��5�2���賮��6��k;�xZ�xý��F�ܩ<\!UMP�����[n��⁻ �5����:TS���� %'����<`�t) 2�`��/��;���?�c">*���%FZ {0̵�4�7� ��K���#�[��wF�5"R�n��~g�v��}ңiQ�U"\�X~�{P[�M�ME&1��M��{���9�id<����ػ��
���|�I=Y2T^���BJ�x=�z����G�B� }�ke��j��xrvy�����3��֌�N�'�,�G�мuf�����}T��Ac���a���+a &��#�ֺJ��d��)q<[.��w���@���X�3�PӼ���#�@�vE�-�"Bfo�����:�Ly]�򕊳O����CncXp��۩�ɵ�ɩ���έ���5��(PD㺻q�mr��=���G�*�WV�]u����obf�8$��Lu��|�!g?�a�'�:+�m��`��)M�R��YC�͵�%��E�ޠ�L������-6���Q��&��,s�)>�Z�+��3����$�E�����'�Rm��&Uc��ތ�]zx�Kh��e�7dQ]����(�䚜N>�����Ix�48�7G>*R�O���t`�^�6c� ��1m�?nImؘBi�P�X��>�ڛP����M��S���ǅZ*~��cm�So���Ү8�c��/y(��nT�1Ԯ�j��6�nW۩	𬭡�'v�e��Jx��� 8n&.D�J#,�q&��H�v�VKd���R�Dʛ�Z�����-��]��t����3� 3l���Z����3p��L�
۵���@��[�����oj�~#{���]GͅQ\I�M
5v���N���-1�+�H6�陇�e��(�����O:���+�
V�!���f��b��gN`�U��ڦ�RE�4���h�W�X�2z�LI�'���F��S����?��HWP)vГ�x������k���J�r�-�G)�ilȌ��M��X�$��2�a��@9��\4?��"�����@a9vB
�����@���G�s�?�B�1���#a�L�ᕽ��;Kg��)�Ef���aT	�/�2�q�ϛ�!Ɂu��v���s���uô�2���,�0J����Ωr4Z������t����⨅��b�9�3?`��6Խf�#O�K|�^2�M7Q<$zq�c�)������=��9h�֭*�K&?6��jq"V�D(� ă���fNeζY��U�;V�d#R2m
l����㼎9e�~����b ~6�};�*��ۑ�F9R΃��T,|�4S��s����$�bS�g�TBJZ�.��)ZB�F��~R�UȳNCY\K�ͪ�3J�a�~���*�"�M����c䣉�N���������^��s!�6�c�t��{���?��.����!����o����=r�i3�@k�ʥ��;�8떐@ң�]�6gf��ٹ- �ɠ�H�I����sTh�&TBܨ��<���n�[�J�� �F�)W1�9zF5�/RA��|�6�~��Hh9L��}��ˇN�I��^ַ�U+�&%N�v��1\�T�3G����DSS��e���F#�o��C�za\�?�V�C�ru)f�L��eׯHNP��tӎ����k��}������q7p��/�Re��88�mu��R	vN3�y(`:���3$��8�ޕ�-� �hR����LyW�#���ҏ^0�9���He�+f�Z�kQˆ*���W�!8Q�ű���t�(0p5+Fv�����ۻn\[�9^mb�ܠ}�xP�=�<x� ��b�٪�F�p��~g�Hv~d��#��bMXn��K��ĻTҡ���"�[�aܟ�8��&mQ�H?��	�P�����=?�����ĽQB��Yg`/��`0!���=��[��k��V�T7�'���K�*P!z3�Go3_�tK���$E�?��+i^rg����t7-�.b��B�d�o06��-�L~
�2S}��N`�U��g(F��L�����;��<��M�JG:���T��<f���jg�m�l,�Z�Ѕm�[��v�p�b<7���M����� ��+-6Y�@{�$��&����b��#��G��{rEPF�}Q�8�"��>	�?��
�-:k[�����4ྶnO);n���Wܺ�xsK�Z�@�k;F-͕J�		.�u]�&�����Y� �C<�dɈy��p��`-L�kt�nXt>g�Q&U͞g���生(]�= fd�/���w�'mtPfʎ����ĐF%�vʌ�c���\���?�&RR���h�U\�v�c9����ҕ�C~k�Cm�(-�/:������+����� y6�o������y��<�O�T�-�����iW�fH�}(OSs��_#�w��Ѐ5�\Ϫ��J>�Gw�0����R�� �	��?5�N ]� ���nzF�u_U��꽊e
�}��/c�ܷ֥M��ޮ�O���8W��w�`;��ĥ\��UDp���_�/7ʂ�{1�@oק�_�(i����Z��k��k#��x�B�`���|;�� ��� �<�i�)S�ۼ7Y �P�5��;X��Kj%���&fa�IN�!��Ȼ�Y�/���־�CI����|"Ym��`|���%D����(��������AO8�����={�[|Bhc�I��I<T�-y~Y�Q�
���7�;�~fh�Ƚ��@!;Տ�ë�_�'2�%dl����6t�H����..��7#y��,B�?s
���·�=�z����X����3� (�)-�Ŏ���bB�j�C@1X��͖Bg�(5q��}�����M�Q�O��S����9���]���s��N�z��=^��R�S�����\�M��γ�#j�1��<�j�]�i ��z݀�*�tW��'u��rѪCL�p�q�!b2���q/�ָ}�]cwv�<x��S9O�R*�5���o/i;����b�E_�:)MT�(l�������ח.ź*�kf�{���1�;�i�%]�P���:��%d��2���=�`\e�눪[���U�е|��k�7�xmГ�[5�B	M����e���K�i$�%�p�e ����*7�f�&h�;KYa�0ۉ�%_��SȎ/��{~���z��<�ݱ��LQQ��PX����X �-�:ʆ��H\u<�֯Wv4��o��$�T����D-�D�)��)�I��w�a�G
�|�S�g��� �22<�o]&�f���͞{����^
��*s���^��t5� �D��dE��:��~�(L���q��Θ�p����pMFYd��
�v3E�����;���a���5��2FB�:)?�j��L����a��kJ>x.ُ�jʟ�������������:@%�W�O�匳t7����ؒ,
#�{{_��`���f�|�n����&�1��(�P�_��ə����+�N�1���6[��nl��� J��=�>��Q��h��|�6	>�ڿ�c.�����bD�ê�L_�����>Q�� �Q.��E))~Ͼh�#p���97|��X��I׻Ս�'�Y�M����:�l�N ��[#�h��4C一{�OD��]g  `7��k��]~Uj`{�\A�������	�������m��d�S~{�F]gMlVd� ���[�WT]��|���ϔ?�2yD?}tpZ���ǋ�����1���p0�w~'�t��o�Z��Cb��%�c:A���7K]eV�ҋ�-�
�J-�\�!��:m/r�B���Z�W~��x�m�`�Vj<���Ln�zX��zf4^��e��E��O{.oNx"���%0���mRzwO��3�N94���>Ke�ա�yE�b�$Q�'a�v��BE�r�a��_�9�L���uu�]����A����K�$��Ѵ?�}��h�-+����c�����
,�T.� ������)k���Lv�{��>���/��%��y����DJ�<%�$]F�p6��E
7��ԅHleת">�(�r��9���&����>(����"^��O��;s��99�;j�[M.P@2�J�C'������Lƴ5>H+�5O�|Q���jc.�֥v-N���ZOW<պ�{�1|l���q�>M�ͼ�qwJ�Z��G���c`�v�'<8�~�2�}�G�z��h�"^��A ��-m�5}��d��v?�-��5������pn��Ÿ[÷�6y=�$�K	�O��5EN���s2{�h���I���K�$�r��nɁ�B"_P�kn��ۨ̔��
_u=�-|T��#�%���2c�SV�:#��x�s��9J='���P�����)����9�>ڎ]�͟On�Ex!X�~D�8f��� C1��P�vE�bBo՝����7�@��1b\Ք�;�!Y(�Fâ;�{<B+�r�zf>�H$����'��X=#��ۧ�Y�G�58������0���߈�^�iHd
J�|�̹�AT��������k黎{.ԑ�݄&���Ҁ%n��rY��Q�@̕g,��QsAůa�D3X�=����o�����LS�_�kVX�jx}��uW�0940F�e�#���:U�G�n����Ey<ӳ�&k���ACB4i֌>�����NN�T#t\��A�#R`7���vE�� @�`�`$*��0W�7P�]V�tF�*&	`�}9;�,jpa�g'�u�R� M�<+Q6�g4A�� $_�e�����iꃬe�	��q�;$�n&�.lRݼ��ɇ��>���ϯO���ʘ�9������ԅ0����F�0dWK\H��+̀���G �O��k5yl'm��7�;�mQh�����lH�a��b԰5��Y ړ��i��.���K���������Z*�-�6�T�~�b@���{��g:EW��qse�}P
�:��rd;�a��R��#)�6�5�-V^	,_�9�O�a+2ꋛ`��Ր����܃�&Y�f��@AC��bo�I����
�>�J6����@P�� EE&aTo�Y�������jlv(�6�WZנtG�	��q�xer�����"LB܉q�u�H|�-�t���"{1�М��;�@�T��vJ��?�z ��s)�!X��L*r��R�{5�89>:>a6'�[z.�w��Ѓ~�r��z#ʾ����q}�ٜk���(�fW�}����������>������b�H���lB>�����˥��}1��d� �&Z�TT� �BQ۵y
��8\���3�-���6&id�F��Y�%�L񴦸Ԍ�@�-z��넘h3��{���-B3Lk�~3���D,�3�>����銪O�q �Nw���.��8��bS8��@�� %��D���]�����CD�8)�������v��>�9�0L��#�(��H_JB	U�w�^N4��H����E$᎟�k�0c��gV�~3l*�?Fv3���:��wC��Ŗ��	�Rq����'�N�RU�Aڞ����ېC2/n�7-m�^�\�ߩ|덌��<��W���^���˴�h�_s���Y�j��+�����R��BZ���my{9E����[���bq9O��~�#l�&=�+^����ه�R�oA�qݍg+�$P�(��^{C��٤��p@NH��Xۑ��儫�T�6^��ʃ���,��Y��m��r�\�R��پ 5�W8�2��k�B|:fϻ��yn�F��������������U��h������K\�l�;g�;��w�
{| b�z��(BBu�ߚ�3H��@3~F9":�+�6#�^G`�h�>�.�ˁ� �=b7�=�Z� ����\�$��3�Zԡ��	s�_B�-�);�'�iq�<������� ��"��VD(Q�X���;k��T&|f�����E�28��0:48�]��w�g��GX���Ѭ�6h��ܻx	^�UHY�>��g,���PUzu�<�B��5]�'�Mbi(���Б�$�m/u@y���V�;<�0S-P!D�p!1O"�]V������ğ�R��I�^H��.���w��î��ׇ�W�)T_J)�[�h]̾��W��=99w����1�b��"�!9���,��/dQ,����h�>�F�#���jǋĉ����8E�[T߸	�,V��NY��(ow�����T4�K��aC,R󶷥�2q`���sȓ�� D���Y�81�ɗ
J{[Ȩpp����;B}�-�g~*d�pm���4��ꭠ�QR�Ʈf����ܑ�I��(/�;g*��I�8pAaFC�b�Rq��B��vŃ�;}��М2DP_���Z�H�.C/�i
�'eu�z��t0����Ef���<�:Oy\êV������p�V�8�/"��1x#U2:R�wɄҒ�[������P�;�ւ�2�C�,�80~��m���V�E	����q�ǜ-�c��tqGD�3Ur	�}��RJ�Йn�HK��ڰsMU���@���E������t�d��7?9���(�/�s0���&D�(NU-Sp� �˓������A:8�S�:?�l��D�rrAZ�Ղ�` eP�a�%2!4�1SB�T:��݈#��80p|_f�A�\V/�O��lA���c,xT���BXS
��~�Rd��W�)Ԃ�#�]Y�#0_dL�mj��+�;�Pz{�I���
�`�:��j�y
��n���SÖ "5Y����w�´�ٹ�6ץ�H��R��MmVhX���d����F���K�ܣE�~ι�G���z��cT��7�q��sZ���}9�ʊ�!m�o�'ּC��ܪ��ea�YqEϤ>�n��v���!��LOk�--._H���5U�|D� ��������y?���/��E��!1y6z��=����62��lv1�ח�����h�����2>Xل������-/�� 6���!�Ģ��^&Uh_^�;I\����g����0�ܮ*��|PKӰ���2�/�Ik�{�$^]���gL5(�в!j��:  r��3��W=�+5�#¬B��f�Ѯ�5�n����Mi0r�L�B��mQX��W���z��h�Hl⍸��7QK�o%&��3���	v�X�佉��[��J\�=���w��&\���<��<�o5��=��8��c8���Yb��������j��W�!A4l��D��[�	�$��{�l!P�_ݶ�\ug.��;�����O|�@�(:��oK���GM�룠eљ�x��x)h}��H����}(��Hz��R%:v��0*
�o�ͥ�sl�+�X^����0o����L[��U���Ng?9��Z���s�Ʀ���xT���ŗXL��4���5�x�ih]�֎����%���įҐ,�U��|��GT�*^!K4�m�D�a��iք�1�����LeK�*q�7D�CB���vx��޶�r�:L¾M�L���0�R 6�����I��ДbU��J�S�����-^��"�k@@��m��������`�zS)C믾jPL"uc�<��\-FSc�Ro�Y`�%�7t��/��������X ��
�|ŭ��T��?����3c.ݯs?��O:�M�ۊj4`I�hT3g�� iC˖{��x`6h�5P�ה�U��Y��s<�0�R%o=���Q�Jx�8K��ʿD�:>>=�q]�U��-
�~�^Rn�����ըi-��5g,�9c5ӎy��33ɑ0��ӏ����"H�Ih�B�XgN`>tc����vu�f	_Һ�&�1
�վ�'zG��Z�N�3�Ɣ�4�{r0�A��r�ɂK��n/zkD&���9�wP��������>���t�Õde�Me$)�lFfJ�u��pN'�ԙ��p�V��b��r�&Ԥ��j�(3p\}TJ�MI�HP91��*q,��0.�yO�b�#p��߳��H��w�"m�\�v1?'^i|gb�����/��p�|�v8���<���>� am�Kpܳ��d2�^���&�r�mI�:Ь����\��K�P��Jg-��I��������q`�z� ��H@��o��FϷz �é��~*��01�vm�mD�l�%����Z�`&\y�Ы'�D@��b�bU$���&1���5�PH�$�iP涤慕���w'���l���|԰K��6q���>����^�R�5���rΕ1VI�У,����(�'�&ě�����"�֝�
k:�_+��Q��7iN��C�ʼR�I�'���,�$�xD)����:�d~��ߜ�]����0��5%:C!x�����1�`�@�6�͒.����͹���h��2�.��ej���<H*l��߱���?�%y��� 巷���LF�K���J^�X| �Rʸ��H1Fa�k]�.1
����e�_��DV�
H�.'M��@,�Eʱ��*lգ�|���q򇉦���
I�-�{22(	ß�&)ۓ�2�^���E��3;�j�1�]!�d4�n.9���]�H��
��g5.�G�E�[���:�P�N��s4�4�$�k��@��<���GwC쨢���4�4�Ocԑ��ȵ������
����-��%�αO���[]ͥ��7co�$�s�(;�ᵫt����n���Y]'�$��>)�˕0b ��|0W�j�ZX4ӟ�}��Gh��z��t��k^H� �������l��A�	[���<����Ww��qk=@��T���K�����"�Ki`��K�OD<����Sur�������Y�����qŮ���b';~����O����P����I)��e�Z��ߺ�WPe�����T�kܥ�0e(�;�y�m^'�;O����ؾt��"X����2@G���]���VXo�r4��*�x񸁈�o`�Dy�Q���;�mw{��^RHa��G'�y5���F
 ;꼰<z�*~���,Ч���4/��½m��f�S�Ï/z ��p�s�ʧ$Y ��v���1pn��_�B��B�ñ�ḩѱ�l�O�8-�)���_@')�MxX@$��l�I�,FR}�}1���ex�1��c5��G�����]Z0��f�7�3����i����[x~T�n9��u%}l�����.�g�+�� �P�3�����)������<��D����-�%楂\g.��o�Ts����$���V%�G�ȀY�
�X6��0���܉�@GXe��W�
��({�RŠi�����a��U9IEO	a�E�E���G���fН�Ut-q�8ֿ[�۽N	�����߽�B驪wPJ�֍��C4�[�I��
�� �&@���n,T�M�tNnui�����AS�����mITE�R��������!�?����1p/Q h�v�I"=����1|� �fgd�o)U,%�)�\�V����d�ɳ���HB����'z6�2u$��c�%]Ȝ{�q�b�V{Y��z�4ucPP��|��B,����솎K�⠹Ђh�2��rc5��Dx�&��pT�$�3%�'Aq��B��S;�`��!�	�J׳.�@�JV��ό�w���߮�^�$q�3�SsiQ����/(_Vѹ�1&Ͼ=�]F.r�=Mp��(*��u ~�8IÓ���̪K�f��~�m*����K�<��h�j�.��Ĥi��6�&,�C�宛j�_+%�<���XC$�)�u�}"P�9��G�>�GA��i|ƃ�֥�ؚ[�����̡����CM�pEm�xp��ǭ�AvK�:�pȸ����YSE�o_$ R��ZP�X�H*Svo�ʈ��b�#�LW<�Kf}���0|�|�w�l٣�.���<����N�Aq�`�| U��-�M'EP��j���Oy/��V7|k%`��rl!�j��FX���P��W�_�H���9�H|jImd�TY�Y��f�٥�6	� �n`zw	���$�������>kr 
�
�	U�Ch��^*f�w��N�%{pYOC������\�{ľ=��D�=B����n����$qo3��M լ[�����J��Vx[IX9�M\-@0f@�,�yWw����$jӴg�gZ d!l�`�������a�c�ki����$2�AD$��\FbDc�iB#�4Rfk���G+5!�azE��f��Vr��3�zJ�V�-���.(t��Q��Y/W�-yӦ��0%7��A[�Y�=������p%*qB�#��N)8*ei���{k�j�3'�]�A�(�Bx����s@��:�#(�F��
=��uh�=�SהTS}

���t+�k_�*ՙ��U��R�mp�i���,q�v�t�I" :A�g�������[M[2�:[9P+n�6ft>0�ל��V��#H\�\t8�j���ly���n
��U7����9��2ƪ����67 ��o@����ﲦÿ���zr)��v�n� &��Dh�)u�6�"�&�m-XE�K�j�	�n;`Pk�(}�&��a�Q=7� ��̞� O_���;]�"`M8��X� �j���ǳڎAC A�e �z��'�<��`fd��ӭb�ث�pw��H��E^�I��|�SӚ��؏�,g{`����|j��V��8Sp��I�y���y���>�(����+����'�_O��%��@R(�=m��Lu�F{�@�3v�zS�2���̭lw��nBk���5�pB�U0���`��?˘�nHn���,��6�7�g����K	�Y�eiJ����Ґj�n�$1-�i��屳G��q\Q��C$F��bD��#c��,���v�R�O��p�����Da�v!%A��j#Z^���/\��bi��*뙲�N����v3��۝F�^׮���H�;�h3-?���	i�'�")�а;���C�V{?Xp�	w���-������r?�s'��y�Qy��5�w����>�͚	5R���ZAx�{#V0�S�P�bD���uѻ�o��
�A�`z0�GI�` |�o�� ���CCH�?�����������K~�y0��w`Ր��	��;���{��U��� :*�Dާ����n��۠��~��k��Q��1��k)�emֽ�\�Lɭ%G����<�><���=��f�hI�3��V�����c������B��EZq����tסHU��(� 2}C�('ѓ�#�I$��k���B���6Dk�7�����fLyȶSO�+�V�OB�����yk�_El�Ɗv\ 7,{e=��o��ʛ��'ǒzrr��A���<�fh���	K�u�U|<�{����}�Z��� 
!'��]�Z��t?�\Tu����U��t����h.}���P��N���S�P�b�ΐ�pS���-��Q���S����ǭ"�b.�JO%Ow;�p�O��^x$������ˠC���*�2�Ϛᢡ͇����Z�2"q�ʈ|�$z84xcp�b��pMa�h�.�!bl؄b��8�µr��/E�3�B��Դ YihQ�/g������bOh�N6��݀Z\�t�'޳�kU�Tk���lڔ�2�}�����^��@n\�+s�2�l~9G���dWm
�+b1���#ltUe��.�߈��\[�\�Ό��n��E�Pk�n�֊�i����_�)�����~�J�ϴ?��2�j��YJ�����[��z���)��~��v'ӈ5R<p�ԳTʝ�v��9�2�"(�g"�+�(��4-K��D�=U�� �|�!^�2Q�������#���yɞ�v���Ff�on7��Ï��b��F��#:���3��В����)e� �\S�cD�K��^�>T�"VF����>�XtA+�8�׽��E�}��I'EV�d�J����_���ur1yN�ѵ7�rY���T�z�MW��Q���т�������[p�n�bDIX5p��q�;���9-��FG8a2F�N��;=,�
���n,��'�t��6����4ik͹d��U����Ί���O�p�V�ɤ�<n;�k��� ��
�WoW����EX'�b`VQV9��J�BeH��2YP\\=���:%�&�nEu�eo��J����q�	I�a=MC��,�w�k�T�[��1�2�-y�	f������{���q��+��g!S� ��/&}O��0f2^��S�X�~���֑w��J��V���%W{oM�%�5�H��q��!\�\*�4,�I�"!�g3f[��A�z��*HN��x���Kv{���o���0��{{�����E�m��k��/:��_�d#��}��m5�ګUa_X���
K�g��4e�}F���k�'|�{�_<�����̝�#dU����n~�,�����?���B�e��}=yw䏳��$H��+��}��
	.�lG(��`�j�Q�Ԏ�q�v��t�h���F�E�_�]�ND���$*�1m�Jj��՚e!;*ubvFW�G���g�tȌ�Q�Ծb!�L�JjX�7�E��9d^�q��T}�s�? B�|i:�3�V�0�R|g���K0��ܕ!?����(��_���B
�>+eۡ9�L���-����X�Ηʜ4��'1�I��q���&>�O��/��=�%�u40�ˆ�������K�4�|q�Axt��:��j�W~�r�~�@<����ͦ_` tV��iC���L�
%*���2Myl�L��t�Ke!���~V�rs�wJ'*ޤ�ì>�
�$��,r�n��L�qzƪo���K�
&�*�o=(x3�}���h���A�5�몚��ǚS�!��v�-l��Uh�2�������eA|-�JL ��s(�|ɈN��V�K����1k5���x�Ac�3Z��1���m5����-*���D`%��B�h�&Q�v���F��ezq�8�T��M�u �Sh^�H:I�A �.��AYa�rF����m���%�0�_[bJ 3��J:�W����mJcc��BD�IȲ��k����`Gh�6����C��%S� �����RY�EE1�w����J��E4�]�.T�z���7��tC��N���1K&&CO>�2�fr;�RیHu|(ۈ������ZE�/���YDG�S�H��I�t����mxTW��!\Dv�c�.C-��U��P���KG��]���%|6�jVDew[$�z�����
 �4����Y
D.J�.���f��y�9L��!2�������e���1��(��{�ʮ���E�+��bl�����#���t;?᪂6_)�Ǟ��bbU��^2ֳx���NP�:L�N6L�
G(w3�9wF�
�m�8��yȹ
��� Z���.�>9����Xiǣ��]n�h4ʾK� T�J{Z���_8\�郀�}܇���`Ȱ��[��njr	�T�Ze�Y����n����^\��g6D�2S�oP��bHe=D1�~�PX?s܌�,o*6s�dG�C܅�t�1U�y�nG9��D��T��`�xx'��o��Q~7^@smC�>���F8��v��bu�,iF�%��S���c�K����.(���odVn��T�(�w4bIf�	���P��n��������MЦ ��r�@'�`�=4(�!�8��M�.�h,u��w�O��bn]�vz�"��*rÁ5K�絑�nL�^|e�l���o��t�j8�7����e��J2�)��I8��m<�"K���!S;���|���FL�>gݤQ"�n�Z%7�E�{�#D��8�%��7�����1�R��J����mw[�&��h,@i��v���g뤋�$q h�
\�e0aBm݁��W���7�%��ܥ��Ď����~У�N�1j 9��u�^��Wk�C�J`O]�@Fy�i�'��Y�rm��t>�嘧��� �vK�E�LK�ɀG��� [�([_�٥A�`�zq�5����̛���w�nz�a���"��N���C����?�;����c)2��_�i �@T7F� �݉�@݀q6` v&�6��)B+HuJ͢���Ple���M3�~���������ڌu�!\�n��Rzf�T½Z�M�B��|�l�u=�Z��@Ι߱ 2K�+�J'�jh>��!���(Tr](�o�M\ɜ(aqBi@kT���G�/>�m[��Z)�[׏ړ�׃�?q�����$Eq4 "G�A��{w��/�E�"҈nD|vѡbVVp�J�2%{�itj�zp%y��/��
�M`Y���8�iႅ���̹����4�^�����џʣnC9�����z���%�K��-�1a�%���%vX�G�Oގ����X���`X��O�B7�cO:�E3P��2~cmw���pe�z�(,J,����������_T��{0�9�*���D�{��f�w ��y� �������\�r���/|�����k/��іw������`�H͚�'���6�������;;|&291o���x�nvkL����K��&`�f3��(>3j��4m'f�����Ioyf�t%87�-�kFOq*56�[�x[���;���>V�T�l�h��g���� 1�p�����z���[���'���Q���6�qG�c��i׹��t�3�M�iwJ��6G���-�35t����X�K�-_� N�3ы��w�M:�=��%�D�!��,3R�mݦ���r<$�֯�,��-tΩ�I:�{Ӂ>r1Y��/���Z���ջ&_I���odKDa��B��O�@I8t��G�e¶m4]rM@is����A��p�U�B8]l����k+yv	�QoX)� _�#fˍ�nk��𦧮�Q�np�u��'3��[���[ӓ��0�|ݝz�z����I��j�������v'%�Hd�	�DF�$R�����r���C6��.��/�$�L���e&-q��ةNA�m@�}�Q��Q�t�	5��Ls��W��S #sK0�E������J#�h��^�E(��\�D��_�������W�!�
��y#�-�w�OwyXp���2" F�π���0[0����mA���
A��G��Q�1��O���濇pz0isy��d������-�	q�Fg��i~�ެ&��$~��m�=Ц�]����,�����1�#KH��=:�<����n?E��ɳ;B�/����Q���v}��G���Z#����G�^ω���I8u�l}faZ��N?�Va�m6�;��S��E0	Klk����y��c�AB�rl�Η�ϥ�R�=���/'beޔ}�{ �A�]%^tY��x<�e�D�CKa9�rS��jh�U�X�a����'�w@M�����x.���-;�u�>�-�}��o��f5۫$/I�����C�!%z���ٽh4,ϓ�A�@l�9�����UZ�\=��8�>Hd���/����H����s-9+n/�Mr}Y�g�s��m���c��۶��n~zg�^)����>�Ӌ.����m��,sv�.[�-�o0H�w����yܻ���scM��&�"E}�@r�FmwQ(r ��fr52f�!��}���!u��3q��.:���k��V;0�h�)ݥ9�����C"k�ƿN�o[ᐷV26�D�!�@�0�� Ok|�����߹��j�'Dኼ�/�z�lx	;٪����)ڛ�iw'w���W�mBW�r��&a�֛I�x��j�����^�D�g2vw�=��!�V�}�@	v����ظ(٣R$�=,]����HQ��zm���#hV���]j��4��{y��I��M��:�h ��kVc��>�gyWT�5����<l���\��k�#x��	uQ��yp�9�D���+� Z���I����ߛ�X+�Q:�c�,�'^��;$^���@nA��_�hma�t����P�t��`���l�y��!-@�ڼ���(vR�4߀n��L)S�jh�g��%|�nh(M��=1p���Ul���/���=J;>
6��E��� 葜i|�=�f�6x���O��d�`�y�Np��,f
y*S_}��,iK0Y|;���h=��N�� ��O��$�?�t��@'�n~����jQ��?Uf����qD%�$�;���J垐R�C�^�dON6>����+6a�@��e|����<�^ 8S���1Fq1)*�N�&����p����_
*I�r�P7R�-��-�茤��(�� �%i4�8�"I�K�)VN��]��5^R�C�W���k3��#�f����!��Q*����Ɔ���D�E�r߹��k9i���),��K�$_���N��V^����p�#`��N���В�˷$��m��W��ב�N;��auz�پ0�#���wsq�O�pW�����w��p�-C��T��N�`-����GIXC�0uy����_�]
�
���8�̾�Z�
�m>Y��-������.k�n�/��jTT=�a��ŉ�BcKr��C/g���;TI=�ԧAO���� �4�d�:"�5���S�0�	��yk�}B�j�����@VƋ��Өl:����	�ef֘��#xƳe�~ue3�vp�����=ꦗ6ȓWA)�^��������6^��ߤv��A��a\��0n7��<�����B�x�iu#��9�QS�x���$������!��`�v+&gU�UV.��fCc��ٛȬ�i@as��`�<�F����!]и�Uɜ���eh�͈.�U�/�8�;YŕD��^�v��L�>������W�+-e�ҏ��/$pc1��sU�V���w"��4����9Z��s�v������I욤͞:�k��S�69�(�3{��J����|�����zn�Wz�����&kh���J�3����y�%�Ŕ�� F��a�s.�Z��~*�<�W�߁�v,�'�db&9�]���I8�N�z]�l�b�!ݒ�F�7�Gc�+̘��?@�MgQ�2շ ��+���x��#Cg݁W���o��E[��R{#/-$J�]Sz%�̤�5 a��~X���P5�L}��� h���b>%�`�]K%� �G99e�j���3�6�#�bއ��a+�׷�FبT�$��V�\����f^��,{d� w�����
N3�9�7�����-#�ǢQ��D�	6��tp�_Eٲ���Ew�X␘�~��h��UU�"��%�>}�$l`�ˉċ����\C�wi��1�����M�cL�ؼ1�o�i�9�E`WQ���-�I�����&V�sK�K�{;y>ػ��ޮ��sZ��ٸ�T�'���Z>����svR�U8Q�y���j���$ob�^oM;6��,������H���ۭr[�}������ɴ�H>i�o-���U�
�{����U�fd�Ji����ئ�����T��Or�|�.��(�����"��tէz�N�)m2=�` |mQ �LA���$� ����U��_<�*������K�!���O5.8�$=�L�R�{�y�eW������$��"@�#�@�IGa���C�|Q���`y�\����p,��=X%�_yx_:a�]��@H��Fǉ�N6LqLf��MR�$6���1���}ǒ��~���+���#ɳ��h�-�;�"߳�����y�	�`��W��̡��ә�����s�E5 ���v{��)4��O�"2g62oV�8�Qۏ���z��cf���ᰧ'�U��r�����E�	1��)�ل��=�	�~�Ǵ`gK�]�?�bE��J=�Աھ��;�>�C�o�F�B�@�~�j��2�4��v���-<M)�nrip?eh�L��ų�c��n�����u�b&x��f�64ǐK�OB��|�m�h
��(W_��������
��m���B�ImD�S� �T)�x�(��2qc��Ǜ�d���H)'��,�?�k��{ܛѳ!9M�P�Fm�Xn�j�K]�- C����_�@@n�������-�;��{�x�P���7��B��b�w/�Z}sg����>�w�T��o�:�
Ƙ^�ɠ��z���(5��J�7��k���a��(��L�H0H�L4$`���vm: ���D��U��a��&�^�}8!?>�Ȗ?�F�X"��>��n�9A��
�#�t�8#�����d؂yj$�>�N���������l�%����2NM�V��0%/cIn%j�s�LvVM��X��'�(q�����V��-��(�p���p�?��0��:�3�������&m��1������,d�a�[7���͸@+(<�R�V�ڈ�����=��qA en{�(?jv��O�b|-�>Q�}�ZӺ�u���
�F8��M4̜=3��w^��1'�Alu�,8|���
���R�1)0���~m��e�l��/~I��
�����K+�Mi�~���U9
�6��?i9���!f�����ӝw�En�����k�ׂ�?��o@����>����dbo_|*�� x���ֱ$������}�Kk�Z�¹&ۆh�����4�9�ԟ����I\��s��-(�$�>���9�P�p�z\�ݭ���3�C�T�8N_�8_���Ҙ�c�\M\)�=�#��G�?����ɒ�~���I�?�bO_x]ߋ(0�/K� n,�NoNK�/��i9ӱ�z��L�i��T4p_˅ �zBGk��ZT��z�)��0wW���w���wF��{M�P��[ۿ�Kb�*���+;ܓ��~�@���;؀���o	C��V��u��c�ϫ�>2��P� ~*�s>�֑S9��4$�2q�qe�� ����t��u�P`�T� ��M��^1Վ�Ԩ�S�IM��0*v��"G檵�#�8��w��n��j���/i��P���-�w��獚>vW��ݮnc��z=�����FeHs��D��N�?��i�h��F26��z�N�
��V5I�ȡ<�ӎiO���D��d��)��"�ڤ;�3= ���s~6�B&N�~탛��Jhm=H��7a�9�H/q��L �)��b"FS"x�K���v�d�^�;��e\yh��VL�[m(�t���,����g�O墅	4$��fS�T��Hqt���/��p��>1��p��)�����[�5\e�8��䥒�N\	ه2MD6Cd�?撍X$�W��.��$\�X��Z�j20��Q��-{�8}�Y��>���58�j�ߢ�Hb��^y��0|����VJE��PX�u�wY]�7m��3Q��U�嶰\5��)�:7;s^AqxQ�!�DG�ڿ�{.�4n��Ү����"_7Նĺ�V�ͳmTu����l���:lȵ�ug��b�ƥ�n�~��QA���">K���AU=A����ܙ���O�Lm��_��7��Q�H@��I/�g]۝K`�"���e5�Ɨ�d!��`R�B����y�[���p#g�\�5.xQ; C�6��L I#�t�K ��)���.h��,������m��!z��w�Y<�s:Q`^�D�x���.?��X`������9_��O�cg e��f�����˞6�#�<��rVC>7ѻ��U�؞yׁ�����)�υ������P�Q�к����x�B:���J\�ۧ�o�����.����s���g֎�S��:/=����m�_x��?�6��a�YI^��,��/�^�8-�R�3dEs:9�,x���fu$�A�+i����]n����q��zЈ��Y/b�_d�HKe�lgT�8=b�O[�cag�-�u�cr
�*�G���Ե
Sl!Y�y����+�_��S1���~j-�B���V���N(���b��hW��!FM����wE�<��Te���\�'�Fq���2���j�4Kcw��)�D��_@=<P�G��5-�:}�E��u��q�Ch�G:���!mh�^�tqW��.��K����"�^x>5�oc���Fo?�GLk~B�\��Y�l<�*Ս.�������7h;��.d�6�eC�VGU����활yx�)r�~���%��"�|�F�5��a����Oq1λ���xMr!��)l`xKj�CT��<,B������1�c���5t��\��O�cKN�c!�� �g�� �g�����{���:[L�]���Uǖѩ�Mg}pvD{�|��FmFN�ғ�f�I�a�ϙ��$R!6�)uT�?u��Oy�j���ii̢f9s1z�sP�|$qv���w̰A���0eb�kX��[w�[�T+$���-�H�1��m��h���CJ�����l��Ī�1���G�f7U|V}#"D�{�k�/s%��sB��~�thz����p9\�L@Q�H�N;[��d��Ƽ�xYW�����:��^�<�:~S�;2c�����2c�D���ŷn�ڂH�!��s�fT��馃���_T� �i4�
��(l���aŠO��;!��J3�.ݸ*s���bѮ�Xb,e�u�Ģ<��A����"������4VY2&r���Tۈ��tz��Y%�<\�
��G]�k���K^Q�t}��R���W�zM9[o����)�;�a�8��Þy�. \t�㻤w���gڪ]�oe�z�{���q|���>�-��{ ����
����p�Z��z`'���;>�빨�M>�9��F�L���|SC��o��i8�=.#�yZ5>`��ɘq��_jb�~,L�,P� ���zK�h���y��,#z��c�=#W�G��� ŭs	I���Ha�iiRFKE7���kI���#z�,ٵ��0a��HѤ_��p��1��>�A�7�J>���y�t��IP"#A��^�yYn�h�]�%��������W�T��[��U��Ү�V~������~��5�F=�o��)Z���Q�iI�
�^�q�R��z?��Ev7pi,�;m#�Ѫ�0��}��q�:�%��IRV_��!���8�z��'�����>���%Vi�9+�FWm��FkDL�!;�'4��H!�}J�g<t�62S�3�w�O9� b��|�'� �^��2Ӿ��3Fao�TP�exQ~`� <�)+G�1���j�g��<�8k�xbZ�j���R:T����J���̲[��h"����r��U&���A�s�8@���K#�1�J�v¾2�y�����[]^��2����
����c̫��@��!7̛�+oiI��T�!q�2��lE`�u�"8�Z�&:Y�R��s�7~d(���\���C*��j-Ʈ_A�fަF�-Y���5��4��gw�0�O�'�ɺ�"�*��9��Q{t|�����֞uJ�4wz��ga�T�*kc$r�;B������Խ o3xq�N�+��*H1b�6�e���.W��
z[���+��ы��:���
:��36�5�d�2��V�)��}l3mGkTA���ڪ����FB����r^x*c���>���&�l0�H�"��e��')��2�!"ϗK���ǔ�WB3�iZ�[n�c=\1k^��
a�mz;e��"2���Ȋ/�X�%ce��I`�:)'�M�ಛ�o��V'��-�\s�����c�<̟ ��a��V��_��Rs	�9�_�4��8 ��k�;Y�\g�9q�Hn���ry��.�GE��Խ�n�K������YF�K�P
6P��<&I�l�c���j��dZ|���'D���?�T-��Nk�8:	1�V�L#�O�WB��_6RY�t�XE}���إ�i�b�kc!Lʅ߭��Q�b9�.����'`���>���I�@?g_�b�<hQ[k�Ԝ���;A>q�@�����x��,j9��<Op� M����i΋t��gؿeJ'�އwz?��¥�A��˯_BrY=�4R�����`�+k#j�
��g�l�C��f�棛�F��ӪG9ye��C|� ����R�p2-RT�!oq�`#�rK��S�J�K*:����K�،$R9m<W>�V×�V�,�u�h$$���ݼjz����VoT.��J�y>:�3��g��<��
����9lcyIG�WA]x�-���$��*k̂��}���� YP�g�=��9�,�U���'FǛ�McZ��x��W��d�ֽ��j� ����r����g���.���C �ML�@����n�v��|���_�L�f��ݕ�C��`�D�\�'����(�s4��P�[}.E�($��C�P3XҀ�$xB�����ݲ�H#F��M��򸹣��Bt a*n�4}k�4NE��{�>����o�m��x$�}���M�{@�	�[̺n��&_�3�Q�%��3�Gt�Z��GsV
V(��zz�e|Jt�P�]�+-�m��N��2�2<�ٲN��Vl��9��fB/�!�"ع��Ú.�(i��8��˜�BO�. �#g���\I��&��T����@^<BW2�e�P�&��A=��6�����`|!�k!�fF��I��({sۓ����������0|��76��!+뚡]��}��!x2�\E뢑9��GzL��˯0-'B��J��s� �(��S���L#�@��f*ϯ�>-d�㆗»��>���^=9-��e$�v&Dk�	�,�հ��wK�B��U2d�	3���v"5�uz��D���N]Z��!��+��z0���ʰJ�G�p�L3��� u���)T�i�8��u��KR�C⍄��9����s[I���~�7��{�_��	j�{�4����@cS���!��>����\�vpF��A�T�0�A`�@0�4i�jI�4ba�Z�r����rl���Ȋu���f�frt�ҍ�⾴�ysr��bdh��Pl�xv��jfe��ֻU1��q6�TI~�!r�YJ�Ӆ���]i<K���m�������:4e�q~�4�'���B��ܔyS���e��BG�Ҩ�ep,��SJ�����F�ʤ���]+<��
���ɎU�4Eou�`�~��s�9��ٯ�/����`��$��ct`	����I���V�p�|u�:�w�(��z�LC{�]~Wu�a�~#F�(��D\�;
�a�DVHQ'Y�,����JO� ���Ӥ��(�\�J|>�?r�drv�?��R�[cһ�Mh�6=��x�y��`�\�FRa���y��G����JF+\:���B�of�q�V������N)`�$r�� �� �A�S�"1��́���}P��nI�6�0�,:߂�=�)�m[1��b�@���c�2[WY�*.Y�d2�>����d$�[�dF�s2��e E���5���#��b%��/'<�{݊ჷ��^J�13D��[�W�VҲ����ａ��k`f�x�5���{C:а�(d��II��3>�o�! [�籍9={NH(ŖRF�x�z�5��߿e��Q�␸��c��r2���������:ų�hs�	�mq1�"Z��"w뽾'v��	ł��Q4d���
l�dB�s�ӌs��Q��Ʒ���݌F������?���qle����Z%Ux�UA\�`�S���7��*��x���>�利���f��r���1\v�.;57a�́�]���|4v��R�,��'����M��{�w�F��&�۷�a��-(�$���,-�Ъ�hC�J�<b��*�ok�����5��c���QH���m�?���7�|]��`]:��o��{�Z�;�H�*��E�D���������ewT�t�H�\�a���瀚3憞\ D=>�✅B�`��]�)0X�ݾ����;O�x�Ys�_��{pe�K�L�B��m[
���N ���=O;`؟!_�=�̮�� /i|]� ��B����ۉ�o=,/qZ�]��1V�w2=0���Q bq><�ɷ��t��7j\��E�s2:���6�ˍaڻ��ObIi��J�;+N�S���h`oD�P����*�Q������G=nL�M�Y�������q�[�,~[GK3��v?�F�Ȩ��y_�Sy�hQ'�AbD6>t���Q�M�;Tb�,v��͘� �VUݣ3�i�cج��?�Pٺp癜�&��"懽����i��Bꧥ'��X���z��2Θ�Mב��}�@~�;��p�Z3���>�!�^2
K����1A$8��.+�r$7&�Mo=���!��@T`s$^��1�_�<M���u����C��{|t=�A?���&�%�lrw������f�8HC�s�w�"�"c|+��8���;[)@.�hb��5�l���
�z��v�7��^AS��_naJE�2�*����#7w��H�K���S��9�����]'�X�7�Q�Z�F��P�>��� �u:.��������w!x�W�~��d)�^零9�� 9og��	^\�D�u@qZ��2?��ŉI�ps�QH�hd�e��g`XKx��+�@ r�H03��� ��d�&VP���Gd)���x�c���v0�زdjoD��mG�0=��ތ���I�@B>HG�<��TN�ZZ�I�B��T�y�3	#;.�ѱ8�\��͂�w�GB������e�����i8,u��!)�\��ae7x��^H�x�!�y1Z��W2�M�����[��z�r'��^UI9H�
a��j
����2A3�bT�w�P��[�-:�fߗ-d�ӝ�ѭ�&�xI������(�ML(a�B�Аo�� ���0��x`Q5�B�(F́���1d��G�b�Yj�AkDk�~���3)	��A�bJ4�:~�q!��5��,A����+,r��\�s4��7�ZP�O�}>�� ��t���eyK���%�M�_/����G-d�#gي�}���lxѧ�S߲ޝ��̹|n{���1�(A~:��~����b�K������W�{ 4�n��4^�֡n~�o�U�n�9�e��q�)�6���q��
��2��}��$�;��$=9y��q�s)zj�JY5��:�f�����.s�6�8o�~�������哪	d�`��z�����X�ssǢY�*�C�cYsȜ�ǆ�L��R���0��;�J�eC��wk�g�H
l�ˍ�3�qzH�ݾ� UHBH|�a�*����`��s���&��냿Wf��{ 3��+��Yw��A���WT۬>%�ų�q�$�q�F���m�0o>+�ഏ�s<lx ����q�r�#��o>gH~�H,S�A@�?.��6O)������_QdK�f�-:�gh�m50���z���n���:	��Gz�K� eљ�����?i��^�+�υ��t`ƥ8��76�ȶ�ڬ e�VMe�>;+4r�?2R�fS�
�O+�w����$�A��w�H�ݪ	�Z���WE�_�����e��!`���S��i8�< ~�h_����6�|'�~�Yl�iza<�Z?n�wg�j}���O%����+z#�8A�G�W/���,�Zq�'� ��M�
�w+ ���x��B
z^�T�AY��v� �91I����|x���N��)��"�C��fc�O����ǡ�L���t��Lj�DH_��������*�Zs�K�L��`�?��f>�k�����t�C4�{?MBKR��v{�'mh��v��"!d|=�ʏf�Pi����ؕG�ȹ~������'ビN�G��UL�6�e�:~�l�GP�"��&��dH�Y9���؋��Ww-�TXp�����s�m��jf�Gڨ�)�(��W!��1!�~��4X��B��?�4H6�&O�Ù��������,QwHQ�M��?��_i�L�r��_��M��k�%����I��ۤj����LY��B�~�a�����	A�W���wa��4,b�vK&b	�U�1e½����]f�s_��_!�Ɂ�˄W��|��}���H�n�.��FW��� �l3'ϱSohԿ�~^~"6a�`(cw.�r��}��6�k�a|� ?-���/@t�WM�9�w���4�R�s�
��cNۦ�B0�_h�X�����Y�j7�u=�C�^�s��t��x���i�g7�T�.s����� Gc?���0����ث ��L8��Y��6���$��>�7��|����(6��l@��4*�*��κ٭���C��(Y�c�p;j֕ɦ�(��Z�݄����d�w+�7��_�Kl��k���6H�DC%^NS��,��1Pњjz���ZQ�o�6)zɮ�Q�����]��lg������#�|��Lv�ɺ��27��n�������-�q �K��Lu��׀���f!���\_�]�H� ��_�8k�x]|�K�a��EH��U�l���.d���ޣp�v���Q�>�$僪�E4W�-�տ�U?uCɪ\ր�����7�~\�#��E��]g�p*�8���GG� ���Ѫxg:��O�( �E`�M��?�d�M�Jnu0o������z�e?9��y�s�S<<�ȸ�"�������FR���X쏥�p��B�s�X����"enPT�UH8�����*$����{?�E
_g�w�=�7���� ��R��|��v��B"%��h~�?�m���\Z�5�����GH-x�ғ߉���� ��������Eōp�����<AW.\���|�F��3 ��]]?��΋0����*����|�4�#"^�2&��?o�ߴ`��Sٹɫ��_`"�-��wz�H���1�6��Xq?��jY���q�-�����&���?F�@&6��d��M��8r��`�Mq���=���z�v{I?+�匲�ö3����Q��~�vH��4ȴ�������L�~W�>����\(��k)�L�5��@N��oL�j-�E2C�c��;TQ�V���JC�����P�w�H�4���l��Ax�^�ȕ���6k����[ákpNoҚ���?�	~A��\Nj�(�s�C�����p)���|���'�t�,P�v��I���Cp��#�;�_�ɘr�ta��g�H�S s�<"c=�~��4~�9�]��!_�dT��+�l�
h<,�#��,�u���P���ǫ�kXbrjԜh�)���˒��O�7������{��.Z� �:���sw�f����K~��1��e���ra����'��K2�5�ǻ�#�����5m����Β%��R���yZ������n�QDw� ֓ei���9�-}��l7ab���F�֧����,׵En��b�^���k�-|Q��O��\kx�rp�PIF|�h��sl*o��Q{md
�LS�v�����6$e*`�#!I��B8
@���0r��ql���\?��sy�u&��_�lK(�$5�05c�ã��Ի��#��Э��_6������¡]�5��""ifMȬ~lB����.-�D��GHi���z޲�QB�X)+x���b�L�9��S���Ǐ9t��×u�"���ӎ�i[����'"�P'�z��hD|�[�oʮx	o�s5����X�ې��-��-�n�L�������:,ٱ�?Fs��Q?���.H/�<�M6�̿����%�YzB�([61{$��vx�Om'�+V�ש��*���e�_���iv&��"Y�F� ��A�-U5-4/��<�@;��13
<mV�����=�2��³k+'V�(0��Yف|��	���X����-C�i}_������4M� �C�b���I�iT��oS�����,�������������i1`(B�aH9�voGBM5��o��gB��K������=�K졿쟞����j�M���WW�*�Nޒ��
��Z��T�k�S�T°O	4�����o����Z���u�g���~Bh�����)��RX�ѽ�E�H�0�"aؙ�2�\c�¹�lÙ�����<����Y��*�u�i("7�i0ʥR����q�J6�ih/{n1�M���Ҽt�r�ޔ� Ѕ��y�:�^��^�9�|��I�ӯ�L@�7��_� ���/ ��]	L���8{�kKZy� c360V�(��QB
Q��i}DO�K�xy�w<�g%�F�p�~��E��IE�� �m[�%�jB�L ]����A�	��]3�3���Q��3�'J�4~Yc����.[�x&��}��[�������)�����a2(�:�8���,f�M3���%:�܊���\��t�?JVۃAt��d�aseRO���b/�����É�
n�h�w���n�2A��CϽ�2̖��j��	���ܭT�f��G�$����DE�E�`��
���������+��	x��n��9I'1�-�
���b%��7_5�K�a Ozu��f�R�7:�����-��b�ޤT-��A�eAwmb�1���m���D���*��&G`_<��XO`'I/�h�n+���v`y��R�tt���w�T j�Z�-�G��XNY��?�aL�Mʑ��rJ�n�-%�[�Yx����gV ���|Ӄ�@>�#����o�b��+P�����\�l���!�u�gT4�:�����>�>JV"�8�ld�P�C��A�6��}<�&�A�zKѪ��o5����S�"�FQ:ѧ����������g1�B��'����} �:�az��}��H�}���)G��Y����yZY��]���<�g��3`@��B�4�;�@ŞD�N�s:��uU7�|S[�].F߰�G�l֩��k���?�o{���&v���\���G���]P�Q���<���v �~�a*0��<Q��H=$r\m�E'WQ� ���h��_�sN�"��&O����}˥l\������l)��!V�$�aG��QH)>9$^z���J��Uq�.M(���%�gL��o�����]=`QI�0�OH��^�Z���m�Hv�����SUN��3�Q�x�5-�ҝ;�%��nv��\�s���_�
gѷ4bV��O��O\�%-�S�w7��Z��9.���a�c\q=?B}��t(�:���֛aƶ�I �O �������;�����C��m�k��f�q�z!�<�U��QsH�¡�*�ƹ��
������\3�" ���o@�FYL��S:7/�'ꩋ���Vn	#�	�B���
wބ��SƳ��ϻdb���<��u|�r����{m�����мA��R�,\W�䀴�5��+�>�����g&7}.�J���p� 8@��&�'Yޞ��(a�^���p���?�/��J8MpoW��ā��g��ƫ�M��X�H���O�:�S��<�y]�Ϻ��m)w�OS��������	J�ׯ��b�0�o�F�w~e��J.�Bc��� OxQ�U�#�� �]�[k�����l�-�!����<M#N]P��%�ܞ��.��/&U{#�m;�f�5x��8��/�T�5������b���HV��>�P���|�S���S����>G>Z7���MVޓ��4¾��4��]/�D$�cE�����ƺ��<:f'/�suU�۽� &���g {���lM�4h�J��RK��$}��ڙ����4�l�3�C'U��}���J��bG���:g��>șgR�ΤZܢc����-����ķp��浚$"/,X��:���%��Yd~�E�>��)�v����v:�t�o��!�9�M����=p9G��} ��ȶ
�E���\G��kIw���8���LI4�@���`��#�F�2��w��կU���Qa+.�a��5^G/cTS�f$*<Dy�`�j�� ���C\X�~������y��/�t_�X�:%�����%r".HW�RG\T9�y~�R��qNEexO�'��x�T9������,��&54�sؔ���5�h1h���;��D`�x�����b1��9��H�d^����$ �,� ��b;�?�Ua�k����,sF���1Rs�7�'�&�����viݕ��7�b
P� 8L��^��%�UH��Yǭ8Rxݍ��5�&��"y���=�v[_Qg�__����D���q�n
L���e!�P�p@7ܚ�ٻ�:m�aNj&q֕ U�R�O�&�ŋiq����/ )��{�V���"���g6CMU������OyI�0�\�����B%��`s��Ť�º��_���K�/,�]��
^��̺4�/���C��#��ט|м��J$!���钷8�6�I�h�~XRB�(k��j�+f�d�%e�ow�����m�Oo"1�.G�*�
�]�""�g"k<���1�P�'�it=��T�d��Ve)���D���|^3�ߡw/I>B���P-+@�WtNP�J:o�)T3�"R(&���vR�D��
��@)�.��8Rí����"��Ǎ�����41n���>�mg�����Qm;�c|��x�N�6[�*@��� ��)��.i���A�|�+ȶf��M@��)ۢu ?d���!$"�2%���c��s)�Wd:���R0x�v\�ȱ��]�G���o��>A�6c��󴓗9�I��L>��bw,�̛l�R�~�hg��� �sJ�%��؏bs1�v�cBw~0�, ���p}F��9����pZ� ���b8���Կ����j��n�]�Tc��"���ٮ������|3�ų_W�mZ��BVI0��qԴD�-��,I�i���`�_�n�
�-Zj�3#�&?8Z��֫{�]�$�Dp����+f���0]�/_��^���H�Sg�
5A�E��G�R7C:ܤe;q3ܿ�x�X�S�hc�`G嬪sKS���|(� �v<u�E������ŉ�m�Q ���a��J�T�%Ƭ�����1GE��?�iF�oUu�%�:h��"�
h�.~R`�T�KK�c���b�1kb���Q��*���4��H�:�]w�η-��5LY��U}\�V����<�]̌�1i�p��s�h1CпaÆ���i���6�ԭ\�vܫ�e���!ˣ-���|2/�<Ӵۊxԑّ��NB�>@������@�-��_�R���Ӈ�~ɍ���7E�Ҙ0�t�����r�e�\�%U���?�u�B���i�H���>MW���w}��k��A�'B�?#Ac�l��ɬ�� �A�%/VzҦǝ"Ou���J�����Ų�ɍzF���G�a;��0��.����	1���t"�X�! '*��+q����>��`KGu]O(���+Ssy�$E{dM���뭨�]Wk�;!�
�c���!�@�����k��5q�0SW��z��N$<%Q�$���3�&�߄��e�t7p��D�q�v-̞����Wr����1K����
�������cH����vm+���%�>�O]�yjMR�6��--��~~���G4�MSzǨHbƓ̈́��8śz�6���������~�����ˑQ$	�/a[H��qT�طə�=��NoPm�!�G�VH�Ȏ{%�@m��gF��<,-��y���N�R�	�Uk�3�U"�K8���!���Ԅ��7c���u�W�`�A��=�!^���*��a�����
N��\�V$3���O���>���KH�x]o�gqՁ�i�f������7�����/E`f�v��0W�s�ыTl��s��֙����A�I�#O�$?�{l�T�D�Pb��pb|.�����iH��;l�cn�M�L"�ΩP ��R=�$� �����ѭ׾�&�A���G�1՗P`m���L����R�g3jL��S�ּN�F�]�A�G�D�NZ�uؼ���b~99�b�8,xpf^M.Ȓ"NG%|����KV�mW�����u�/��mZ���`6��;�;�Q�a�c��U�
�aBJ�ô��mNB*�usN�fS�$xu��᱒���������J��W5�z�x�6Yί�F�S^��$E��.��ϐ��ئMG	+d�z� ��U����Ӌ�[(TB�)����F5�4��QN�R��ݴ�mJ# smI���w� �)O�6�T����?����tyxj�U������W�뼢D���5dm��]��@���������ԭq�S��Z�?�o	(r�?��ny>�۩k��������g�P}�l���Yu�{o��F�G�."�5��p!
������_�é�M��]�+luQ��ʿ�Gi�0 �D�'���G;�a,xfj3(F�B27�j�y����p�z�#�&�I&&o��۸�3�Z ��x]NF��q�z�VC�a���5�|�!($/]@+>�HLo�>V�p:�;,n�K���2�_=�WwDr�����#ݡ�SR��OY��B���7U٪�25��L� ʯ���v��fᙂ�Y3Z��@�=/f_g.j��q�w@E���?�ī����g�th�<X�.�WO鐬�O)��5Gv���5}r��F����^���>~�;���Ot5����!��[�4����K2�_�܌MAd6o>$�i��`����;��u��>��!q�=�Z���V�5am���1�b=_�T��I���?���i�1��z(�>���Q�M�86�?@оy�q�KC	H�WD &]�����Pi�1A&��9�M�7�$R�Ԓ4��WV�Y���h}vq�$:�D�K��?A11��Oݏޚ͏Bg��f�Chp�-͟N�M���n��_�3[�[����mr��Ց��opp��'�N>�Ϫ�����uD���\�s��<������p`���*k25�uN�X�������Lnf,I�'��]Rs��,�gX3�H5/SN�ၔ��MΆ������z
bI�<��S��������[Ԡ���4��c2�>�v7Rqk��b�Uu%������g,e#�^�Vr�b�}#vO��<��}��Tf��߭�e��𣗳r ��}B��f`����͉}YU�j�ܒJ|gM��I5K7p���I=R��Ǳ񉸇fO1�@Jt�J�GI���d���V�r�Q�ʥ�Q�	�T�+�m�E5��u�U/��C	6�s�~ ?�i��3�"-�iM3g9`��!�CdO
��3�	�1q������5��=׵�},�?�ovH��Br�7)�$���%?L��̻x$��Lc1se(�^Xߜ��9:} �kC��id��m
͞(��h��#����d��UI�J�?����:�%���<��f�-����ä��)�ӛ��"fv��C������f�]�%Y�:�"0Q�F����t��jF��x�t�^Rxa�U��ڗ���ց�h:����a��O4��T>�@Mn����OW7��@�>��[|v[�B���=_��jXΥˤL�8t�{|oHR	nD��F| � vY�xt�q��e���H>�v�p�+J:<;Z8x#��N�����.g:.�ܸ��L�'��!�<�2���s/�i1P+C��6!o�dY{,q������&bi�|~�)��%]v97��
���>����Wa�>�?��P�+z9�LH�！5��&��Q�<UX74���C3O�J(��:C��d6�(;?�~- �V�sV�m��˕�âĺu7�<>>�bn�+'iᗴE)��$�ѭH���y�;{D٦-�<�܂`紳���qn����B$��d}a��PRh��p�$��z�Q���bݘ��4�us�~�ޓ�u�{_����,��Fȕc����u9T+B��x�gI���f��G7��S�Y�(�EF���}�t���~AI�8o�ʲѬ�������6���yy3����հ�`@N(V�}���t��� ��>�YP�5wd҇���B���^0�\�y^B��̅�2{�t�	���jd��ϲr ]�	�+%����))A�:����O �԰c���Qt�7�K�x�>��7ڏ
 �ߟ'����UY��͉���B-��);�y�zX�h*j��W帤�])��,bqϠ�
`�8���D�B6@����0!�wyR��#�� Im��a4z!_�b��?is���;8��� ��?^�sO�?(��79/���fr3��z�,c��\O_%�6OB����J^�G��^1�6
į��'�3�����x���U����x��E�O>�4<�n�Wvqi�g���t����=,6ٵ��D��D�7����0g�u��0]+o�����z�s��e�C8��J�����T;q����ܹ�5	��Ue�Q�|���~iP��I���[뛄^�7���d4޼cty3䰀ʹ�O�|�~ �בב�Hӱ�H֒L���I�x�*X�����ϑ@mp�Ny,޼�ς=m��h�02�tDX �hT:y�%F�%ߩC�6���P��$/���N=��+���,F+	j*^�mn�8�n%ٻ�<:L�l�{�=��<�_Z&g~&n7�%��I�
�ǳ�Q��l��VP��c��(r{�W��A}򼖿�5E��bO�l�����B>rCz�"��V#��q�i%�CD_�{���*�(�b w q}q�@`1F!e�=��t3��-�
ƈKYtP����܉��������Ɲ ,IrS��YM&D�2���G���rbG3~���6��^������RD�:�*U�</�a7��:�_��:��T����y��#=�r!D_��Y�NM��v3����U���2��n_h���<C��_��4�8Kʒ��ژA�T���N	s��d4����=���/%���?UCT�ɦ�-��k�a�:Z�7���@P^��z���E���"��� >7��M�q������Si�h�R���:��<0�pJ��� ���ss�1�0ˀq�2�j�vd�ܕ$�� ��Q }Y9p��/��Y����\�
=�{�������l����;���d/UY�-٫��ŅOW?��FkD�*�h��<�a�Bu��Zy#n����3I����Y=l��G(lU�v�E�ax�F0L��2��?�9��Ҧu��R�rFw��\o�t�Q�`�cWD�0z���x;���kS�_|�Bƨ蠛C��w8�r�ίk"��!Q�Kue��DC:�/���:jL���I�]�a:j.q�zf�
�QL�ZRE��3v�Z�N�**�u�zP�nv��^�@Z�N`���pZ�yP���c�|^��N0.��x �2��� >HmAj+aygk��^z-Qu���Q�6�6E �H �EX�2��'�T�j!�.6�ݡLՏ.����뚠Ӗ��`d(f&/>�4�6Ϟ�D�]����5�y��4�e�/��O��d�F�\f�$`p�wM�⹪� ��+bqƳ/e�y)��E��|�������xl�зs~��PO���L=���}�o	����q}�`��cu���y�����kb�{������0�K�n���C�3b�b&p�;��TMM���d��x�����*L���*E�Z�:���'����Ը������ ������-�L߯`�1���ݮ�ؚ˪Sۆ(�=�^'�V^i��S�7*��6h/�j��ǩ�x|k��qks\<�̍4��πWoz*�Ɵ���s2����7\�'8�EZ9n-�<Q(EM��>����TRƈ��$�V�j���o#�3����d�}w�Zr��C'�M���s�5�!�[���A��&�D)1�d��-v&��Sv�r��t�Vk����J���4�j����^�+��_0_���"#6�sS@����f������5°ۑ� ��
>̨m�ħ�c��+:�<��D?س��	��nsd��g=����e��q�^�M�RT�$��Ue�`��.�zPnTc��X䤂��8��|!%�����1×g��v;-��\�4\���T��j��ٿP�\�d!I(�^;dmt(����I������;z���,�f=�ndvz꠨#����sK~B�N��C���Chf��-��C-�V��Jx�YP��DǶ3o�Y�*����e��B_<�I�%`��K�}m�-��c�;(�乒Fj��_�A��/��y���9>.��K����Bdy��H�4X������2q���l�.֖ӊ�M��ȹ��ͭ����zh��cu�^ps�_E�/`�S;y`���΁�}v����h"|^�����3n6)./+�j�o���϶��Fͫ6�2MmC�q�ي¸A�|-s#�#m�GL&<�\ l,�!��^L�^���g����ÿx�.�Zݿ1�s�Ŧ���nuqs�qU#���I,T�N��q*!?����=G���Ą9W"�ЉLT7~�K<��`�\��B7v]]�$��Be'>6&�|�( �	y��6�-���榑/4K��\�Z�k	���9�f�/�ϛOoVI�G=�[9(!;N��Tť�4y�L*���ف�C�Rb à��ެ��tB?�#Ʃ��}8ՏJ�z;�I��-Qk���ĩ�f��q�KTp�5/�d庽ޡ�z��g��]D��Q�a�5񅜨�qym�v㸉�/�o�`9Ly[����F�f{�Ɏ���r�`�=t#�pY�� :�GR4;��_����o�h��nJ8�7�w�Q��O��pd��+/��*�H\f���t���No7�s�έP�r���"'g�z��x�-���=I�����Ҽ��y9P�~�}�P�����*-����0���q�_���5ݭ*h5�PV�����xx����̙`�����b~�4̶�	"����N�aO-t���p(9x)�^�U�n#��?b�?L����2�0*T���D��6�	�f�)g��Թ]��t��Ѩߤj9����S9��VMx����g�͠���,���˭Z]��r��$ӉiT��� p���zHVe���a���mBf_kX
.�fɁP)�-O#�����Y"҉�	@a���E�g��/����.�ҽ{r%�eI���+�
c���.���St��"���aUO����j+$/1B����$pI9�3��d)�Xey�G.�)�u����T���T"/���j�˓nݻ�}қ�ο6�_W�":�oz鲬��H�s2�
V���Ӡ�Z�}���ʹgo�Xp��7Bn͛��w��n���4��,K}�3EVbc�� �s�|����6���?yȫNr�SZ__�K}�)&e�A�LE��|X`2�T�,�=ì=����H۫��*�"��R�H� E�_vW���i�=�+|Nh��/9k˟##�+\\���(�a�̷�Ʀ�T&��cS��c.u����o�@�\-}»?l1��︅U��M-FY�5�/�4]jޠN@V����*_�@7M8�fk�]);m�K�.�i�3R�#���Rue���t1�)�����H�ؠ���-��VD��rx�I.��~�ki�~
�����a���v,cJpY���J�̗�/�T�ᦢ|# �e���[Jw+n�`�[?�o��.�ڴ�TGP�h|	�>vYG���߶�"=�����Pm�j�,(^�Μ�.���`9.[L[���B@eiؑYvw9��1��<D0R]�`y��rB*�r1�b)����P�
�ϳ��=���@��������P�����to>e��_zRA�͵��̹7�m/���
�찶�l���0�o7�C�J"�ZE9pV�6�
n��S����:�M}u�`����{I�͔r:��0��J`9�;���/�A:7`{ug3��,ĵ!{-�Μ�w7�	��ܨ+�c�Z�ԕ��R�i�o����"˟qH_��X�g�҃<��Ca�҉RF�;�A)/�53n�w�AV��g��zey��^���@@+��i4E�So�E *�z������`�O��+��}���&}^��ZO��| �t-�,�z�����A�U�:i�d�R;'v���Zpw$���#T��P�C�xr��s"��%�����H��'k;[�����/�g;��mkm�g��U���oj��H%�'�^0��Ɗ�s>~�#�� k�X�^@�1�s�Cv�Z��+]u���rk�>G���_�u(jIf��i��A��������RIG�i��7�B��*�~����iG�d���#��C���/4짅O�S���q;"� �g��Z���(�(�v�$�G���d>��ɻ���ĎYUi��q�f��0�B����
"ܩE5#a����!��T�K,��Y.9$�j��J�f�n��O���/��|��`e4���f�U6S�7i�.�B��i؜ZU"i�}F5��"��s��<[T� �o�}��A�K�`y���={�Z������j�O3�t�]�O�?<VԹ;�`�(�%�
���UT����}2Tt��qtl[x�����OQY���co�U�O�J�4t9��/1?��h,V�֕��T-U�p�Z�o:88�ʊt�R�\1�"YOȰ��bY�/F�\㍵.�=�5[�ZK��ܸo�;������'�0��⌅- GR5��9���i��S+O�g}EMl;�oߞ��S:)<��:V����9� �1�Y�G#�
'� �H�޽�̠��d�����_�'�mݸj�*�*��G�;�3��{O`���tg.wJ�Z<�rqD�G5p����	��g8�Z�r�ջ:�Rn�S�<������>�)�9�,]
(dD��J��qr�Nۈ�-�3�M�ڞ��/<d�2�{�( �¾KuD]c�b�x ��	�wY��<��f�+N(������dbO_��#�gB*x�z!��_���F�t+��E�T-o��i"��e��sY �n߱��ʾV|P�m���Gx����h��.c][�)�iP���"����[�Z����Y)��ɸ��
���Zw���x�^e#���3�I<
#��qH�����|״i�F�h��(��;�|Q'�s�д�aeȶ�f�JH�g�ID��f�t�4�8 {��d1X�H�|
n9������Vh�]|[��2�+����P�����<�(F�Jt�Hƻ��r@n�bHUu��y
��N�F)�Ѐ�J^�MC{�#\�d��E����-�����'{��ĕ?��)�-D@�w����<AKn��֙�����Z���ޟaN�w6����a_#���1�|¥��Z8D/���?:�.Oq!Ј=�KU���;��� ��� ������nV�?[ڠ�}>��+�5�-<�#��'�cF)0����hxv6��G�u˖GA̐��]uj��*�Rދ3��|��v���s�#ۢ�u߷����fm��u���GUR"��-N�L!l֫�vg+�Na��~��5D�����ë���]�x���ԁk�j?�Fh��l����{;�u�XBORy�s�jR�Uc��)��_4u�ՠ&8Z:�G�9���jc5^E���+��hjFx�K,2Z��t
��̏�M��l-wC4j�0�[hb���U6�DLG\a�խ=g72ll�	d��6-���Tn� ��N�@����̱��)�IE.�E�Ӓ�_D��^NV~}��חZ�|SrR�@�H(H��	�����JN�{�r�)j]\7���3��e�8&�-�+`��I��G_\v��^�ζ<U�=~�Ysk�k}	@S	Y�ؓZ�d�^�"�:�m	����:��B��[䘧Il���t/��CN�6QΒp�2:��� f�^i�<�ԛ�b�CΑ4_8 ��k/	i�A\)f�w��V:�0�Sa_I��V���n㘗���>�Z�ґO���2W�]N���\c}�H*`;.��	�6�r;����Q m��l�Zt�M�V��`��>�A���/1�~���)��#hl�ƃ'�$,F��SO9SD^F*.�2ꄥ��	���հ�����G3�6��ye�ÿTU����o����@C$�w ��n�����mf;-u�Q���1G�V �G��ZCU$3[�ƨd��?[��k$��h�w���+�A^�
ϐ���maT+$�G�a|�h�N�B����Pf�X ���_�_�o��6]�?z5#�����I��%]���n6�(�&;��L^��;������QL#�h.��7��>Z���ם�S��r�����s>:����>Zaɑ��t@�/����B4�(�U�h+�=�(8y��;�[�~�s�mΝ ��C���AiNc�_�,�V�v]~;�"+�d�Y��k9�P�g����'=<F&[��c��GP%0�S�HOP�֏U��%7��\�$��d��7���)[� �l�6�0�MvB;NaXZ��¢��<�Gs��ؠcj�`*I�YR�P�b��<��M�����N
���R5�&�~�|Yl^<ma�R�/>$��y�i�O'�ђ̆��=�A��a�蝆���)F<�4�T���b�[A}�D����)1���WJ#����!����m*<�nR�F�f&��P���fb�o��)"��g�ꧠK�䪑CK�
��.3Pk������*���Z �M�[^a�m���r�����0�n�3���[��+��͵�Hz1��%�
_F�O��({����M?��IiKO�r�Lv~h��R�<�馃	��6�n(ε3�����,��S�f�Z��~5
��lV�^Fi���S�v�v��[t����G~w���_������B�mLBs��P
�,�Dk���Y�(nz�� �V�kX�g��,�-��d��(8K��O�G���2+�2k�ݟ3������%�-�g`I�W�sB���2��g���.!xڄ2����8C�.gM������׾lgi2��!��QF=j�_��N����nce��5�뭆(W�u�m��`�T����IR��M�u[�S��U�,j��Vÿ��W�Q��ä>���F� 8��59�p;ր����n6�qSc#(~RF#��$�ݪ�I�|���E�8{T�7E3�^��tٙ�'� ����AתJ��)�r��&�ٚܣ$���z�H	��u(c�=�e��so�vaqEV���:&�;��c�3r=J���5�腺71��r�����K£�Se�V�;��\ϯӏ�̓1�\ʤ���)'��e5�ג&��C�����)*����.���us(k��I�e�+�#?����!��Th�'����n�wi�q�/ ;���+�o��5(j�x<V0C�/��Ko�-%�}�/wr��L�{GE`K-2��&�)�����oy�DL~��&	ed7���x��/|�͟�Z���Q��-^��R��ٰ�1��|6���z�ⴰ8H0�+;��R>oK�g|�2�n�
��C��ڷ�؁7cDx�0�&��r���]��,'9��e��XLd��T(��K3s��/�$��'#(�c&m7��շl+�"��7h��8^�U1�`��K=��j~h��-+Tf�u�2��_�k��O �^J-^���0u7��K�9i�^����7F�q�+A4�'�c�n���`���7������L�GT��LS����~'���H�+�H��9ǳq�RX<2:����*���dj�Y�^*�m�Dd[�"V}i�vYJ���xd�� �h��V^5k�k�>�>,��9��r.���#�R?K8"=��W�0�+Y�'������b)\x<�?��{��{�����܉7���C��œD�� �f$�a��)�C��\K��f���~�W���$�A�����i�;��D:�84ۊW[��G��bͮ�����O�yS+��|xc4~j6�v��b��	�AP;dS)EH�X3�]y�N�S9Q�H��[R?*�/��?f��<�;���27t�p�vd ����������P��vCk����\��ƥ����o�]�� Z1���+{ψO6UP��2�u�K��;XEx�[�x�T@�� 3�3��T�;��+�w��g&T6��"*D�������E ��+}���ti�-sY��ؿ/Bt	��,&T@���M�T` ���z$�
qW�8RӨK�j�\J��C-�7lX��iM �����[�6�����G�$�Y{�J�H/�GP.r����&!��*���
�-�;���`||󆖬+����R��3h\�9{���ݭ8T;<��,'�׏f�A�)ڣ8P���5�72��4}�5;T��;��r��&�Т�vN 4X;�/ӳ��6+)�hM1de����.(z�(g ��O���̍�p��$Iu_p%�\��z	K�f�(��$lHV��ӹj�@�PZ����c«��<�0FmX�\����~��B�G����i�i���������ڕKS�!3{E��"sE�7y ZG����Cǌ���?��[��`+C�3�(-�-<�UK!w`��.z�m)��&-8ո>J�hgT �Y*��gǐ\+f1獉)Z��ĉ��A?��=a��Sg[�t�@%*�$�&�l�����G���1�yk���hF5�_�@N�Զou?O l=�!,��%�rJ�����2��b\I.aKB�2WcDmܪ�j�dVȬi�w%� �T�Ah�GM�+�R:���F�#T���t5��L/��RA�*' �XTX�}�A��{˲j�&0�v�0Kl*�&Z��]H��\�$�J_�����.��;= f��K���'Y`��IG�������Xp�_a[��ؿ�M5�Ě��)��Mw�=��u\�D����i���� F|��L�h��ۜi�^���ra$*�s'~y�;b#�!S�Y"�.9�`ju��,���&(?�H��0*<�:Hzݴ/z@8j���j�;bF��pܹ��Ɂ[Pe@��cX��MH���Ic\s���!�ׇ���4�Y1������5�F@:���8�z����ݪդ8F��>��C�rǬ�Ň#��[(l�'�f�������M�xHcO�}����"���X}��
_�K$+r�
 �-���K��`�:�/]����'2��ٽJ��)�9�n��0ym	�7A�:&/
4�p���r�@0�ҩ�t.>�f,	L�=�2��V�c�z����Fz�\���{3-6?��ו��4�;��_]�:�N}�"�yѣEF"o¹��4���.� �B�S�e(G��q�au�n!��C�Z��NǤ�c���r�a=8���6�81}���2^Q�ߏ��0���{��r!�Lֹ��W����͵�KV �T.`�!"��������e��L*V�����i]��-ُ��t o���wU5��s``�d�N�a@�%�s�����ܙ%w���i���?i�^U�&��6����^;V����y2�=���󪒲<�`�� !b.bY2ާ����P�H^)�qz�P3L��B1Y-J���}jB.���l1��6�eɕ��	G�L��vX�`��Ȱ��h��QA�:�#��ً��}m��۫�
���:�kȘ���:�+qg4�
�~֫6��H�}�C�|]'1^��R��C@������GL�qP{A#�]�e�/Ξ�WJo�;�^n�i݃�e�ig��o,����ɿ$�	�yS�ڝS����M�κ�b�ΨX:�nk<`��Z�a��\DtY���kCU3�wK����i��Z���rϴ`OUp�'�-H�\p�3��>��lp˛9z�k�%�K8�J�B�j1&�[q��`GU�5��KIP��}T��E����+;�4}b��̥�>�E�MXyAz �#.����yQ%�rBV�$��m(����C���$v`�Hw���*��W�}%3�fo
 5� �K	\����G��%���+�C�HJ�ԚTM��?�4[|�*(}��B0]�N���}j���/�^�)J7�%�!l�^N�c�q�v_<b6����|xl���SU�v�P�.����Y��٣2�63��S��N%�i���ԇF)a� u��U�1U��&�a�b�ٞ�g�E�U��#���kʛ��������dM����H�햭��� ����� �16P�]��l��{E�)��;�
X�x �����Gﶽh�Y9�.���g�s��v��]�n�^m3s��b��;	y� �P��K(��_y���(��#L�����݇y�Ĩ'���u��R��WYV�5L��ͷ��b/�X�	t~ob/��ti9J)��7ğ��
�B�^�I���J��Q�e,c��)�`tjUr����$��|��B��Ҟ�s�e*FY%J���zF(��u^t�n��a�m�K^&�ޝ�Q�u������10ied�|����������_{>5O�������^L؆sq�F��esrGZ���4X��i`�(�S�6v�`�Ė��mFu��n�Z��A$�5��|���@u�i玖z-�|t=�e2���>u���񘉡������7�G`{�s������.Hn�Cef���&��}/�lA����<�7q@� _.��i�[��:O�JP�g�
����i��ث�3��L��Lt0�SoKt��+�°�a=7`V�(�=�ȸ4+l��8���f�p��n���`|Ziΰw�Aa����L���/��#_N�8ꈢ��t�?���x��I�:[�n�SBf���� /��ٞ�}�.k',�	2"/�{���O��8�m�=�������Zoԛ���݀G�/ŀ|���w�шa/7uVsw�?ucs������ˀ�"��c�~��3}��Š�7-�0U�@���U|P�N�k�ςu3����Փ��}���vk�([����(���0��7�1"N"�3���q|��V)92�kZc�7Z���Q ̖�� �X��鐋�)�g�QO=�|x�Z�(~I�-�.e�V��#���~3́O7D�ɀ觃�#�e�s#���?����*7�>�W�p�f �^�>��������Mq2���d8$�j�eLs&�Y;�]~U�:�
�j@��t�3И�Hv��.��o�dyb �]X���d�A��?��+��R�5�.򪣡���t�~���V�ti��nPf�@�9�*X%�$*�4�'N��	i(�Y�?�Y���R�./#�}�A�^`s��)\�榣h��;����<�=G�>�	8/u�bo�{R5%��ۓF�	�T?��qă]b�X0CٟsI*��S��w.c�h&����)w�mGSD>�Q���+W����"��&}B�C��s�.D~�2Ę���o�%o^�|w#����r��oo]�:7�&�e2�UCk�.��5�O�:�F�(_N���Ac����1��J������p᱊iLm�>�a���K��y�|$�Y=��.�HC�����B=<ʦl{Z�,��8"M�ߪ���i��kl6�a�.F�!�*������(�R�������Mwwΰy�2�ucPJC�����"��k��|h%ȗNPB|����Ȁ�:�8�F]�|�U�X�k�8�9���������ͱj�F�����pm:� �q��q������o��/ߧ�k���5����Eh�+����Ӎ�Z�P�M���t����|ˑwXQ�$t�Q�+{�As\0IVf	6���ֵX�^�غTc����6�E?.�$}�{����������?X,c��\��#��ֽ�d\�Tj��2^��9J�;Ֆ=���e������	s=��Ǿ6���Zm�b�]Y�z����2�E�r�1�RN�cMO��i]a"6sC:�&��~�}g��ڛ����V�s�D	~6ҧ5PM��xy�U����}���	�Z�
H���ϻ H2W⎒熘eU)��@)�bu����!`g^An��ф����3J�Y�u'J�F�v0��� L��g�,��o;=+�}�'!���|��Z��cJ��p%�x��$眳��s� c�����6�_����Ճ����D1�����*�R�f@(pj�?��/��ؤ�������WSe������5�}*�!A<��֗���F�(*z�]O>·qO���Ѣ�����&�/&��W�t`M-�A����\_�̲6{�2�]9�ݵĦ��c!P�|Tƃ��@�`�kJ+ۮ�$����F@'�|p�Ev)�e� �
�-Yq���YF�V��R4x;C Jl�!��g��3N���O�g)e&�q�P�4(���A�k�늈Cȝ��ϔ5�g\�P�@�SH\,Q� �`��y�ﱛ�eT�q�K+�^_#�uc���'}�'B!���3�w8���;I�T�oey����	A�~B�`sʶX�-T�U�T�Y^���B�ɐSD�Q4:����)0�Ɗ�b���� ؂5�~���g1Vh=/��]�s�|��q��a˩�Q��Σ���˥��N��z��?�t8@�4%G���Ԛ:�K�a��ȑ7�w���Y������;�-���M���|M�n�ѵ�u�Ӈ�V��A���
1W�:�3�QQxd���3���d3�f�
�Z��<��f����)���lC�.yn5౑j����h���c���ؐ��J�(2�*�g9� �Q���̲EGh~�X��:�4�tK+�#���������t�kq���TD��-1!�6MR$7��[2�Ҝ��qU_W��d����h�����}��Z���釭WYm�l���NF��r$KD3hW�H��a�S��2�Z<����v�)@q�Y��|���u�rX���e�J���f�h�p��ND��y�l���D1�\j�G<u7�W�h6c���<Eڬ<�cߣR���R�r�P�q����	pJ:�ø>(�g}wLb$�����^+�'H�Z����.�cF�D-2�w	%{�ʍ|xCpO&T4�e�8c�;�ɦV;�-ҵskVN�,h�s��Xm����XO+��*.��*������*q��&j��8=�{���jƨã`|�)�Ĺ���k0���&)�Rtś�7 ��L_JQ�;Om)�N&w���rJ�Y��!4�����
�G
o�G�?)��׉y��l�!�P�w3<�ڈ&�P�Ng����Զ
�
�Q�����Z��6���|�#ÜO:%�T��1/��co��V&�9����ŔB��
��?:� ~�~�����䤓6�3n��Z7��t�c&~miq���U-0�o�}�������$�V��;1�)-�r;2/��w�_��J_W�Dk�'����7�k�u5>�d�l3�Mer�
 ���Sc��m�@ q�!��q<KS����H
s"�4m ��͐��[�Ĕc|/��}x�&ɥ��⸤�k���69g9�O�,f³� ����@_��9R6���%�0)�"ɔY�J�BWc9?I.b���Dn�*���0��l�2��԰@!������7q��ȹ�V�VK����Yߥ��G$Ɋ�ysb�v�w�&Ɂb�RMJ�������`?�"�R;^���e�iS3cX����]�l��r��Mub��i@�_h{(�r�t�w����w�c�i��v�jb�*=����H�U.[�&�-���@��f�����dnr`9Q\���Hx
:��!�x��ZxZ�
{(�/Ԝ���ɋ�=R��k�8ۏ�/��Eׂ���N6���|�x�@��#F
��rf֢�ޕ����#��L1��Қ���!G��/e;ܯv���$@��:W.+�kޘǎ&B9�Lanɛ0��jA����ĞQ ���X�,^�/��/2�D/�_�w�\a��[���sH},�(�����K.�7�����xD>��z�,�~��#}G�D]��J�0<k�;\F]����q��)ɩ4;�����8+|섰�X}�!����'�j��b Y����\�|��p���c:�ד��!����rs͊k�ר�1]��&lTU�}E�J5*Aޢ���q��Zag�p�`�;rE���F���4�w�_��R.�+�3Nt%i5� {uُW�"��b
b*,X�A��=��������-�� 1fBｹҺ	��j�Sx��Q���;>u�Px*�Q%���c��3��M�n�LTp��Ƞ<�³q�w����X=�q�%�Cn��������̩r
5�`�v����0ϰ��.�������U���v1f�!Q3�/r��t?��̔�=��?zh���Z��=�s<"N�������U�kxG���=�I�OI`;2��@����J0��$��+W%ԭ�K��:y���kM)z��I�N����:�D>�`[�ǎ���������F(����<LQ-i�@{n}�w¼����GJ��� �A��]�v�����-�m?v�s�$|?�~�����p�s��]��L�ң������U�ᅗ�Pjrk�h\ӿO�����0�#��W`p�w���g��z�n��Ԗސ������R!����]��Mi�zJ?_�K����hщ�O�T�F0��6�� m�x����x���3�S
V�����y9cOv[ݼ���g�-U��%L����y>a8	I����-w��5�|Ҿ�
�շx�/M){�ͅ�h�����OL����m������1i��D�����"�&l�>T�a��	RB*	ͼn�9�@S�~�V�OӜ�7Zd6�%|���`��i����]�6n��3���
�O5�5C����|�l���cJb��:,����:C+�]t[�Ј׭���4�c�1&C��оO֬��̦�t�0�jI�58��"9��VB�/�{r���������%��y
��:p�pأ}�듫d�;�]ߐ�;LR��7����r Z�x�����ub�㱸傆���x�6��<&|gݓ7��}!�T�2R�d!�v43�8}�`��U�P ������L�=������GЍ�:e���q�H�!��ŵ�;�1�����,�e>��M���\�-��-lu�^#�Ӳ�*�#��&�)q<��sKm�C��b?ȂF�\��L��]>���P]cDN&y�l��K�=x��(�iW�]b�[��������R-����{�0O���%��p�o|��E葝�i����Ϊ&0�/@Y;���۶BQs�*Ƽ�(=w��rU��f�q䕫��
�>�aE*|kN��:���E���hJF��/F�`:����o" 0yG�`A0́)x]`3��&�Ұ�@�v!�~�,4Oլ�jGs���q3Uɤ�aQ%�"'��T{&4Y�$�����p�Ӫ޷��ҽh��k��m纬�^�_&%�u��|>	E���Lac�܅�h�7����JN
�&��D����mj
؏w�D�x�CD��ٺ�M�"-���~>$��z���h�9��bS_�k��������*5P��Pl#bhĳE^��i���(D�	�1��#��AN��w��*k��N<Q�K3������_ppi��i�i�p �@~*#��1����Tڇt3�i�:3�1X�R��F��N����O1�(��<�+�W��h����)T+���V �TU߬�{����o��avĹ�����U�p�/��u��X��,�3�C���8��@��s�yl�=zL1Z�������]��G��I�j�T4��!������Hq�R��'��U8W��d8�	fm�QQoE��.���/'��Vðf�r׹4�醋ʛm�<�N8��qAi���.)�?ݍ����pch|��,7���,��8���MB�_*��!$�-���e�$�iC� �.QԳ�;��$�,�UU�F�b�@�!V��{���M�?���5����z`�%�ۥC�n��AC�����VZ��7Ob������y
���h�]\LA1�F8�k�a��I$·��N�]��>u0'�O|��`�s�tI�9)��$�Mk�pԌ��X�k�e�������LzW��3�en!b�k�;�KXx�`�G�^����9w����X�۰H��TX��`>�Bv1m��χʿ������Q�  -?/�(�����/Dn���*�s�s|;{��9Թs�EM�s�*�����<�	��~�,S�����߂��d��_$�)Y+ė fP����&#h ���4V�S�5��?���cU�%�P�DN�',T#��*;��f���'^ܟߜW�VU:��Q�Ϯ[�~��Q�+����-��l�k�Rx�`Op�V+\�Wp���`{���n��-�����q�͌��ô����2@�'ՠ�z��)[��ΐ$��J�|m�������iz޿Z�2	%/���`%���aC��5��^.Xr�^K�kX��9����&0�*��G�_��b�n�Ρac�����O����k�ajm6y�6ˊgOd�3Ln=�ϡKЙV5>tj�Q^=Z_�g�rM���kZ�e��^��,[*�Ʉ�'A���+^4�e�~@���υ�.,̺���j�Gs��V�N/-u�ָFq��u}�jAg>���TӢeBI����.%�kǛY-�M]�d�6����m`�e��ŗ��Z��I���P�2��E���p���:|b{	�9�Nt@�	zHr(yݣ�'y^�؎��=�9SHv�����⡱��p�I�$C� �V��3OT#�:o�1��?�lS��Fϼ���������E��Aӥ�N�s�iC�!�B�j��Jn��W$�o��Pʙ�H�k�&�G��2H�"E"�=Ex���[��kiEЦ��׽%���λ�G�P��T|Sl�n�7��U�Ҁ|�����c۵
�A棵�ߙb���:��Fn���]��C���z���wѽL�A x����
�+�X��4��s���U�T�?�������墫�3l�Q�9�g�u�q�t�NNZc�����c�e�Ah�\��)`�f����ZZ#0���C��r I�%p�<�@o/�����T>����K �O ���5!ɗ��:�.c����r���~�����ӏ����~��8�J@艽Q�yߎD���gy�ѧ �B	����������;>ULp�$J���H�mP��5��8����?~;d�xi��2~G���-��q���qL��t�mDYte4'P�ȶm��}������;�HEK�q�wqS]��U�z9�p�E�Ζv+�p��N\&%�)!=���@�����_�C�8dpGwo%��nc�Pp�3r�6�GH4�GO�/�Q��H
F�<� u���~j�1��)�r?"1�$;�+��.�V���0�/&
P~~�����DHK#y�k��
�	��[&_�1�
�y�_s��4.ܨ)�\�O��7y?e=��݉���@���-��M4�w������k�:�-��z����)n�
vo�b5㨊i4������E00N����%.�<��Æ�+�@��P�@D}:���p�5v�[����W�̛MP�f�OId�+�Q��^a˼vX`R�P?�(��ք��U~OL	�=���Ȯ{�N�����CZ��g���΄��q�,�੔^9�TU��g�5GTb�y�hsAΘF�5�����W�e U���7)�N����7!�4���vh���_mm7��Tǰ���I��컇��*��>:����"�Q��t�De,�G�>�����$���qM��v�{��g*�n�$� ~$Y�n/c���c����I�J���D"	L/w[G�:F_W��櫓�;����.�������-�m��:Q���%C`�����^�~�e��0S�e��[5jUC�n��w�ǳ@�?v5M�ǩ�E��'�o����V������ �3�.li�c�n8��V��MQo�ۼTNr��I����j\��Ѡ�x�va�-5�-R`RVH~�{��O�g�8�H��T����5���Q�8~_��:�G����IX͘��j��a��M��G"�yh)HL�_؀����	n%J�����HS_Y����Y1{�5�1~"FnB�yN���
��Q́��s�|�^�Y�ֈ�d����L�Y�o���Cֽ4On N(���oL��F��--EzV�'9���"�V$������l�� ��7(FD�̛��Bf�Z����\���vp�������@>!x�8�	�s�T��tm�O��F�U�w�pr0oJ׳�4���gO���,;堑�O\|]?p�\-��,U�Ґpxl��_�lJ+�/���U!�/Z����
'�b�+���7Ce˲1���/��5@]wm��� i���]��B�Kx�"3�R�w�Y��ᗷ���K������M
R%��*��5�dcx�	o�Q��&Z:�e��j�x����l1)t�i�c��-�b*X>h8��Ä�h	H �9wM�q�'�:t�SF^��a8z�u�D��.'f�e�ө?d�!ؾ�����u%�+j���^�տygV�H��co@R�f�ͬ����/�n��G���~��N��*}r����x	���_��g������J)��<�����_��� ��w�@w ˇ��[�ވ{�`2u)�pD��hw$�P�'���Oky���A�z��#�%�E�c:�F��U2�DX ��z�Ҽق��v��(�7h 3j���y�w����/#�q�+���l��+��fm�`T�f�O_���#�2�6�Θb���=�~�� ��t��Sw��V���kL��M��h�հA_�)4[/%!;��L��[޵��B��
�C�mIk�P_����?��q�v��K��#�#ôv
m?�{-{b�a�,��ܹg�v�B�')���Fj���[AQ���"��ڳ��%�yb�H� ��Me�ֽ,XF���w}=Йu���E0�h� Ys]�37r�^ql����38"u�׆��������0�,���Ma!����..O�3�*REVv�dgۮV���A�<vO��E�2�Wd�|2v�;�����GTʕ��0�6�Ou��e����yJ�@��l���p���E��%E��=�=�Ȇ��v1>YMꍽc=6��?A�/oCⱻ��0�|_�{M1�7_d���4�ݰ4+=]ɽT
�	����[��� �D����H�1O'|��܄	�&?�A̠���%�z���潄9��}�N[��]J�ň<��(i��"���z ��Ym9-`XV��=}UB"y���K��A.���s�-LM]����``>4������=�����d�x;I/$ )�e���1�WAҖI�m��z���*S�+Z3}\.�	��� I�@��wժ�װ;����e����Zg���bm�W^��3h�0������C�9���������_��6�⃥�4���`1��'�<�����!�g08o@=��(n8�^B�ѱ<�8�(4ԍ��'����C�Q�����*��U�ɖdY�5cS�����6�+b�sU2����}jrB�9�wY�x����,9�!aI�~�t�H��*�ȝ"	I�����L�*F��ڦ���{=��
s�E�c��<����R �^�Ξ�m,4�0O�Vuc�Oh���C�U�f��K�Q�X�~�P{iIq��A������usAp8�6��܂g>��x�q�OE�O���.���j�gJ���e�W;�.S��K�%k�̠
��(���O~�:���i�����i�7�+�z%y3�BH�?�5!�/�/���9��y�'HS�4�L�e�݆a�;V����$�>B���v�&�	b}�c�>Ykv,	c~66Ԉ��"kJ�mnx���u��Gˀ^S�2ʦ֝Нa���(ш��/��<��yd�V�nw]B�����
Yfa�^��qכPmL�d�\t�%��,Eܠ�UA�+&s��h!<���:�w�_���zόM�Y?)�5���q�-Ь�0ߎ��
��v������#=���}�fb�!4�H�_j�	�G��tϮ����s��p��.�M]?GJ�����G�u�oݩg�!ҫ�k��JI\�l>zXz���tg�з��eQ�� Z��_�yX��`]������%6�'H2�D�p�Wq��/,*L�=*N�7M}h���}A�:�3�qB�b���T#6!tX�q;������UT~HB�Ēχ/�mkAj��CȜe�Z8J�S'#�q�i6�����\J鯙:='�w�^�E����_�Yȼ���_nV'��v@~��)?�hf��o1pA�d�ģ��(r{�bti��M���ҫ��Q��1���CW�j�ƫ��8� w!~OO�p;x�luN`�N���]F�Q��WD��y-0ም�S�l|BqP��NG�6)'h<�(v[ӄy�+�0O7@��N����Lc���$��qŧ�����j�S#[^F{ǔs`y�}��ba�]G3���Z�<��L}��t�o���祪��?�(�~���:���� �K�*K���E٠>�%	��s����Z�3���T��"��:��$/��#����i��Tz��f�>{�Le�Tݝ�i�-�����ϣ�N�����{?�HX�xCjc��F%��3����C��,�
]R%��{��js-���1��%P`�ڌ�wu��"3�QKɲ叼q���P�5A��񅌗C�@���)�|bX$��ó�e�9��^4�hwa�-�65$#x~/�{[�c�J��5t��=5��zy�C�Qz�C���:OsDvS�Oa�α�.tV<�w��|!@V��|a�nws����k�z��0�L4`�3�	��|N?��a����,��AHi��-�,��t�n�L`+|�{�W���b|���E�fq�Ut3'g�����;8GH���^GKg��<�wJ~��oP��d�'�Z�l���)X`|�%�_F-�j�nS�K�W������q�_|�{����!YuHL/��-dW�ƈ6�o���o''��9���O �=�zP�(J
�� �B���t��s�/�����'� q�ԤƐ���h���'�"��(f���*v`V�\���j���J�/����i�;��HKڀ=��1�.��8�>�8��(��?Idz�,䋷+SaBc�g|�.��L.�xJ�+ѿm��Z��%���z��e9Z>�$N��ݭ\��UŬ��E�H.���Q2٤\�ci������ �d�s,ZN�/��_M�����)�2'�ɿv8F�}�Ta9�oS�Z� J�A�fG�k��K��A_w�8g�,�����.�R"ez\�Q�c��z}���ɟ��HC*m��ӡ��Ō*��;������/��.�S8s.�Ly���vz�tsfrAJR����cY�G ��#_�%Kg'Ԁ�U� MkB=ٱzM��٧���i�f�gV������PĬG�p���LP�=��/�Y<��m��9^��/ɞ�u9�=�;�32�'~��M�!��f��hL2\)����*��BNe�=��ZI5Qfs`��W?��*j)�C�.���O% �W�5c�I�®��M���Rep�K�SıJ����PLl�}b��]��JLإ5><��ÇN,޳�DDsǔ�vx��F����T/6�vh�ߌ�ҏ$�?����C��,��s��k����_�B>6�Q�r��Ԕt9�|7���Zu�N�-�Z�n��N��3��Cs�2W���q'��iU��s��j ���"�����N<>�+{%�؇�o�d�"C�$�����qoG:����'�E��~���Tx�sK�h�4����������vI���E��P�/�	]��.�(��SK�3lٿ�#���� V�R�.��K_��4.!h���য়�@4���?B�EK�$�UҺ���|)�8��)a5�i�A>r�ZiWQ��'�����sħ�f���fl��/zT���s?����3�	�2���~sߵv��!����$9��Q��gF�%O�e��Q��v�l�	��b?�z��g�j6E9�Y�uj��FeW�)�iPq��׸�0�%E�� �]B�����,��k��`���H��\=DR�s9�}$�ms\�t�hR%y�X��ӊ��Y�	z4����µ�������a��N� �2��Z�=GN�kLA�g�����J0�}\���P�bm˛
3���/�/nP�(ǌ�b���ᢷ��u6 �z`�6EaD�Q0�fn��s���j�=7�>Kp��Ŏ�f����:�j!p��*P��}��4��+����t1�'���fM)���b>�f�M���?谒�2d�f�3ٜ�^GIF%(O��(Y�m���E�i��������G$x�kᣕ�lhլa�a �� �^؆^jᒹ�Q��.W�w�/$�*->��|��8��3�!�8W�-t7�1�l�&I�%/�0��;���d�־l���²+��;a�"n��L���7�P�uL��4p'$C��;ok��<7GM����{^\��r�pJ�})���o�	�E�$K�Nx5�?⦷�����x�یM��m��	"��w����H?$�S1�e;9��.T�m8�iUC!ܾ�Qv�H�*�����tIŌ�<Y
�t�ω��K��F���V�>�����S�G�+����y�v`Q���qa���9�bK5.SDl�s���߮��)e��5m�C������'V�������;e�E���b��Ч�A`��L��.$��秚�R7?��$D@|�b����4tm.&�P����F[��a I @Fl�1U�-�5,	x\[�܎�u��&]Ů�?�0?�V�Z������EQ�a��7�^�0�s&��1mǍ����U�FU)J/��bm�L� "lW[�7ЭM[� ��"�j�t�kk_�J�Ͽ������4.,�G�f���h�{RJ�ӻ?��S���Ƶ�<�6Guծ�[��sO�p�NC��$Ir�|�Ä��bn��a']�F���Dp�e�p�x,���t���� wP�^�i=oˣҌ��꿁'GɦKk��y�$��e�i�;�����ϣ���1�}���{*[�	%E�5ug3v�%G�u���h#�j1�Dl�Vz yf�H����Sk֡���i״^��*�P\�+��b!���ԕs�e�.7w'���&jh�V���۽���\�h=�Eָq���ǆ�`r ��d�@��0�8Ia�I�V��b�NB����T�/�� �o�j�-y��9�E�qa��[57�����1pI{�U��k�ut�;h�e��;�M:���/j7	��`f���N}6�l�:��|8�xV-sֱ��ϭ��V�� s��Vi]BNw�a���
-��o۾E�W���R����"���)��;;|KU�Cj����fz�{0�+��R���zg|kp��<�o���)p�%���^�&=h���b~Dە�Y�ח�'�l)Q���{���&�q���t��><�dAt=����O��9��
���֒�f!t��S*ѡQ� F�tɘ��ʦ�1L���n����j�<����Dq���Nקބ����JxW�?y2+�n�4����5h;9VH6.{����x��9;�[��$��lE���߉�$�?��u��G�yI� ��!U-�,�w����A�����f�4Ph?��󑷧���_��h�WR�*R��bȒ�Gtk�ޓ@,�t�o~K@�[�.�ϓ�
H��n9a5����U��s?��)��%?�T��n��UR
˟o��~�eQ2��	͌K�Ӣ`�|���0��D_U�Q��8���� ���|n� ڼ���E�|��Ƈ�$v]�F��x�˥S=v�ܔM���e����t~ܪkV��;�Wz�d��_��I�%�+��+U�zU�E�H,������0-���'���nC=������G� 15���_�@z��Ӣ�8�F�T�._uKCY�q�CJ5�*��ͯ�.H)��������ǭ�BE4�mＳ�� �zMk�z=v�w��K��~7�6ɿ��N.��1�@ KG�w���`]�6���F6n,��4�E��BYk�O��_D�\yr�.�{+�*:eޜ
�A��'N���g����R%�V:�ж��P$,�R/�����Nlz/ec�$�a�iW�k�7��5�-jCM{�i۵K�v�t(�u��|9�� l�R����ND�����ps�J���N�Ҝ�VL��n�̱b��5Vvi�ۘء:sE�z{'y}0nΜ̰f�d�H(X>��|��O�'�$�F��-D�9LA�U��T<w�tF��(�Ο��W:7����.��+�Q�ۯ�]-j�
d6��:���r`�^�0�!��=UR�����=j�V�ܫUv��S��M�o�aV�:C��f�Q$��ZD�j�i=���FR0f����J`n��������P�"�ݚ�e	���HMo!����qb�Ͻ�6Cیu�m��K3��L��Ӆ��t�a���y�ˌ����9-A��/�7��;�=F�!���|I5v��h��|}�rدY�b���C�z�����ŉ�U��PF1?%4xT��������7���o4e�m��H�b��!�_#`	�OO�&�{� M�;C�"���j�N�3�רT��M��+�@�S��T���^�Q�MY����(F9������`�:p�3Bm�F�}*h%�o�pF���A���q�	5��b��t�9�]I�������"!���g)�c�a���*6��6���;��������CZ������|����]I�c�vb��1G�J���c�]>���#CVOZ/�����[���W��\�ǹ$�������i8��u�<AZS&<�� )j��U�B-�[�Y��1q�Xĩ
�K�5;S�=1�dDE������*F�"���׈��e�.rn
\�b��Sr���B �@<�Ո&lZŽ9��x���?8���vm��@|,��b���CH1�琬����x�?���)������2�ʲ���򛧊���=m�<���#4�H��F����lդ���*����8��|����� ?���(�}	��^1},�	~�';/�P0�C&�oxe�!��/�Q���0+#){��U�pX�L%Bm��s�|�s�I�j~7����G�x�ͯR�zp'�@���w�n��`F��E|��J�E������S��O��0,��}+�ο��hִ ���ɿ^~��`���������cP4("����}���+l�h��ᡇ����?t��o���Յ.8p�N]D�o���w��IF�o��yًu�똏������|3�st؞+Q�%�~�>�Z�>��H{f��c�sR�k����d�d��w�*7FE�qZA�%��$�'=��CƻdF=e㜰$����=:���βmISd���VH�Z��T�v�MI��AOc9�j��*F  �%x�n�ܟo��c��P�8QL*+��r�p%��rB�6(�\�o�z����L��T_+�1�+K��&&MM+'�F�&��u��$��*/5�c���$J��v�a�{ĝ P��JH�;t��T]�So]T}��+�r��v�8~5��y���,���9ۧ ��e�_cK�h���������c 2y�EA���ų�j8ޫ��~o-�rZi�e��>'6�"�C/�����Pz]lkƺ�bЃ��y�_�>%�'��J����<tx;�I+�Z2��T7F-h�լ�r'�H\P�0)*X��͈?�#�����C�����,�����
�~��+U�Ac��y�{������fC��\U�LM�v��,m
��K�d�ͺ0SQR��+,Y��<�e�E�U�Ú�Xq��ӗ�, P"�%�qJ�m��SF���*����ћrNh�Q׃r��:@������[���d`����P���AQ�,�#A]�"pZZD��u�'��Jm	#����v�Y����
W����n*ĕ�/T�(k��)�L�F�w�z+���#�X�0:�)k#1Q�׮�'~���&����M���L��m��D�g#�j�@�����/K���϶<g��I)�Kث��u
���lS����h��(��3�uV|l 8��P��N8� V��DհXM�Z�ɑ�jJ�e��9���Ӫ&���a�+���V�l�7�!7�_"�ʆB
�)����?7���*�h,�_��l(��up����&~���=g)c���0~�K#l��DsA�z��"��1�#T�
�����ػ@a���VB��S��dNi�b��]�^b�BEX��Pb!��B��M�1q�7-sX}8zg'�z�&����D�\�Wq3`t��o�`�p�L,U��T&�Z
��!>����k�;"A^:΍���������jX)~��4��$.IgV�;|���N&"|Xz:�ejW��*O�[\�d��<u#�+����ȶ�B�{��ۏ��<�OMJe&.l�:���5I��d!
|%Yҧ�/2�.���Ɔq��^�æP <Wn��J�aYUJ��O��@)r�l2T�����ױ�xK�c�{� ǦQ^�E��7���u}�I�0��ER��|� ����~2N�2p�>>K��F|�'Xk�)Xq��;LFs��S�Hk0���7�z���hR?\#Q����#�q������2G?�W��7�TlǞD8�t��"b/�-��>�^�#��M������|:?Un]�d��k�#a���F-�|huA��S�#��3o#NT��Z�8R�r���"N#��ou��#|;�T���Iek��M>��RB��Q���6�8��8Y����j���8�m�?V35��u�}r���t1<Chl��pQ~�f�e��UqCf�}���exM��%iChgFKu'�1�H�����n^����8n�n#sU�K��k�(ۋ�n��k��L�>��� ��B�ð��Ǣ����[3���_ԑ�zO��Z��8���s��!C�Z#p��vn��59�G �A2�
v̺���P�O\ �B7��Ó�ӊ�+P6�'z�7���l�c�{�a�DT�������EDJߒ����RY��:�4V�
�A=��~�t�A+d�UΨ �)����3/��8�L�nk�4���*�Y�JBm�]���|g���ʤ*Sg9A���DO����}.�����!�֬�6(³���v��-s�bp�l���=/\]JX����5���Y��yb�_���� ?��X!�K&G#�����<*�a�0n�f���"J?~�V�g@c����Q����\ f%�����<�C��0_
�%��{-��g�.�@��4,r�Gˎu�_��Z�߯F�߫SFG��wD��E3f�3eX� �qi��̆C�y�e	z~�^]��Q/��{z�n�exS>�9�B�WuI�>����r�/�1�e�[9�z�cb���ӏ\o�ɄI�ዟ���)8d���y4���tHP$^����/�H���j�Қ�m(�]��^6@��/A�B�.G�t��͹X�Nf�<2u\��_�N���ˏ��η~*�Nf)`qz�͢K�J=���s���Gá��2���OJ�NB��Qk�WԮ�$xgWTzjՁ@ǜ�^�s�9�F��P�v+m\��攮T�h�dR6))ԄjJ�RdYθ�(�T[Y��49�[������t^������<WF'�(���o#��J����Uq-���ؙPF�d%~�p�]!���+}^�dI�X���r�A;Wlx�b�5��(�C�|6BxƴN�G��g*Bx�Z��"�ߕ��y*�(�e>�Q�-���X��m���4�Y5��d�xI�!%����ߟ�c�p���kx*揋���+�ע_��%*�J�u�,�ǌ�X�,��O/��:�50t�#�2��x��Y����=`��J�XE���1n" �J�u��"��6v���7��ư(@�s&�뻟�#�NbW������M��n$
Y��J�+���&	�9�����߼��d���GN����V�\\{ƶ�[u�k"-ʤ'=�\�N�ʻ�i��*���پ��Fe��p-�|1�5�b�+���ԍy�1
�ê����� }Hl@7��t#��46�̝�jr�C��{�ZA�sf�`���bM�57��( �[O�q
ݦ�˷Q��*�C���[�r�g�P�N,o�M�'L��e�q݌G:�*Q0g��+Kܵf*��p���-B�H��u�ĉ^�ե&�xBZL�&I�jv%�*r~�/�&<�%�䫍XCM+=l]cN(�{\���U�&/��U�^�4��)�`�i�U�OAf9�}�h�7��s}ˋ�n�)���5���/��%���O���!�j�E�7����b��&�9�C����>�=4Ȧ(��X:Vl:����S(4�?����ֹ]{�3�RZ�m���0{����U��E���8XZ�jJZP�X�ؐ�:�'��Rz � 0LU�M1��جc�5H{�� 7��@��qw��6K���#��e.ɴŲ����x4���G�Y�Џj9zA�<c_P��hi�
��� �����8�m|����kJ[������o�+6����h6���g_}.����:�2�����]S;y!�����!T�<�v���8�b����'~�"u�fÊK�����L9��~�����bG䯐��~��+��&���8ngv��������+z�_��n�QH�x탙+�=����mm��9��HA�CR��˞�?}�oU���ЮA���!sʟzt������uH�9���P�tc�������<@ƒ���i�P3F���Ê����HN��{���}꼕+�kW�f��)��dq��jYL�
;�feSH9���hV�pE:��T��9�@�����an/�����������ˣW��;BlX��2�V�e���)�쉈i��T*䓚�IV�8+0��t��;�-s�8����	��ӝmɰIĩ���nN��ɰ� l��o��F�'ۨy�:�J*�VYr(��p0z��̅f���g6+��m�X���t34E;mlJ�K�Z�5�]��7�"o���I�pK��v��*��K%HA��Ac��t�H	7Z�w�V[oxr�૱^��{<C���ѡLx���2K�]�/�J.,���P�[��>�W���j�Ȟ]$�p�%���k�o�u��#N(k���-��lb��K� �� ^��f�1z3[Y��uh�
1����c���SӒ�9�A\��2������䒬p��beJw[ק
 i]RR"cqG�������* Q�@�B	�)�[�_Zv� H;�`�vM�p�nn%)�^�H�#����6�
ԗƿ��)]�@OgC5���]DܚP���D[Q�Ȗ<}	Ny.u!�eV�<Q ��9H�b��Ә����s]
#�3挨e�)�P���9gR���Jr��qj���������ir�=p�C6A=p�RGK���Dڎ�;�/C�Ăi"��ٰ���tf��B�J�#�W��(�+(��}U�ݪ��s�Ɩ���∞E��7	ai"��Z-�*T�5xb։g��#jX�m�'��\!,���AW��)�S{L�ԝ�H�V-�'����<ކYP��}+���2�Nm��E�bl Q2m;l�mF$b��ץ��[����>��������<B�԰;�X\ g*T:~g*�!�(�]����������[ND����3b��-O��;��&��ى�4vIY�#R��ʊ�b�{�ɻ�;+uWh�F�s�֟��e�y�4�]�, ��\��6�6#�#�p
 x�R���O��d��C��ǟM�i���0�s�F������t
ܣu��J��O�yk�i�EjN��vs� 9��!	l�BB��H�@����]�Rm"�M�	����Y��@h�c�m����oK�;�5��gb������夭k^��c*����
��F��6pJ� 9�K���a�����@��"���36|�Q:��W��� ,���L�Ī��7ʷM3��4��h�ޝ�z��\�4�}È!��m+��[�'^9���x/����(�r�G�� iWj�1�fX�-4<�������Б�/���:1d�/�~�#���j�V!���T��G#y$�� ��z.��M�ʏ^�!�_��0���.堣��FC��ؔ}~�4,.�� `��������Ky66��\�C(ʳ����ꈽ���7�%�b��h��� ����KR�c�hq�m�V
��/e�5��'A�+��:�X��p�3ȉD<UKßi"P#��R�����3�^�V��_}�Eܾ <.;�:��Q���l�M�� OҢ�A�k�?ۏE'���T�lL4P^ш���H��}���(�������Qt�q�!����V�XP�k m����hc��f��W�
r8c�O{���OZ�t7�_����������\�K���]W��#��O����-յ���m-�ɀ8t9�-\aA�{#`�	]�1J3MHT���[�Rj��p�Û�Ė���V6��e�kjo���5��p�(�1�Ƚ+�PN b��X]�J���HH���t���Y��cw�
�9]�>�Y���@���2R3b�:���*��v#;��N�X���Z��JPv��ȵ�z�@��U!�27�N��,��$?Њ���j�eW���RX5*�[>�DI2p��tP�4�u<׸#���'�|��'���h��I��$@p";����Ho7*_Iv�Xi�� '�z�TR��r�D�����sN�Txf\N&D-��z!�b�{�Vj6
Ea�9u3ˇW���26��Y�t� ��@as[_��?�F�K���3���2�[���KJN_F'����a���p���F�� ��ʞ�	:~�f$�o�w��g3��2�܊q.H�Q�9avr��'�ov��o�,T�y
��0�=��SV��iC�w��ĵ��M��Mu2-����1ُjb@C�j�������2�U*�q�K��SI}+T�M�Z���˳V���Û;zҷ՚���ߧ0�Q��W,��:����B}���wUѾ���h�簗���)������4%�h��K�}���^�M�ħӦ'��OU�KI�gs���C�m��t�d7E2B�����G(�����wL}Gr�ի��vH
�˟��#��w`X���;Ȩ-hHp����r9����"��l�R�qʧ��J��OL%fٚ�ߗx�������_#��W&J���Vwޫښ�1im��Jr&6�JT�Ɇv���}�]ҕ��?]\��E�ށc����&��Y4�����~�U��y��{���9�"B�8֞D�\�pH�X��Na�1�V�Ĺ����/��ܼ�	���,��#�bB4����+��E�
)�j�%<6д
"�n=�~5�l$h��ik!�ᶃ��9j�|�9�����A�j�y���>�J��[Ts�N<M���o�ٻ��+�HD�ڥ�̄���>PC,��j>��%��>� �w����5*��8A ?juW��� ʗ�(�;�v��S[�<�W�2[MU��;1��A��Dc�Ao����{J3�.'g(�������Dߋ9򥘆o���<Q#TC8lK\���Mքhߴ��F���8�n���#d�=���q�>� �;_,�ˋRk�М�m�k jK�p[�/�.�(T�|0���V�+s���F�C���5gP�^��I��Or��K$���PM'��m��U������W�9^4l7!�C��]Z����`%ue�����+�\W����������b��.Ė-�p��W>P�^l�8����xl�6K����vn�6 }��at�\Sy�i�������&j ��u��L�P����lE`����1��js���H$��6�]+�+ч��,ڶ�_�����"�Gx��g�׹��߾q�`�~�?eޖ��N�?������j�p��W���dx��^�J#)!z�uSF:���p����Q�+��0i���q�\i�]��Wݸv���(�����y�֏�C�@]JoL{X��������$�ui���%b��gk�������v�;��^+^;M�e��o�j�T� ��X��-}:#z$`us*[�Н�uP����ŝ�N�_�9�%�7H|P���e��HI$���e፵��+D����c���O�.�v�&Cyi��חo��]��jNVX���6m�x訓��yc� ��.hW�L�:�ZX�S�ʲ^+<E�~��}iۖ�%�ה�c��$���(ذlMLͫ�!�H��+'�-��	����qF+F�N13��qֆA5X�\�������Z����'�ZL�!<kS��(˜J��J9c��ߴ�+�]�3{�O�an����ס_���@�,p�9�,��H�A	�j�ccc�z� �D����
]�ck��_�k(�R1�C���FX٧L���A
>_�>"�&�R��tu?�pN��(�J����DP���������-)�J��GG�)ں�>��J�E'i����~�c��_���}yE#q7�m#���ϕA�)KZ]���IiM���9�@��pV;AN�L� Av!�ӦB���<lT�g��P�BI�|Q�0�	�(}��ƁشA�(��� �8&)4�Uj�����$G�<>~�_��e]�L��TƋ>sA�Z���t؄���E�mNp�+�P`��O�I�I�=��]l��B��_�2'��W��H��ȸT�Z��H�l�n���Q��L���dk��LLTu�<X�@�--lɪ�F�šU��"%d������Krj��M���ýoh4`�e�g�!�dK8�6�h����tgaZڴ�qb��,�}r�d�l�p3�9Ȳ��6߄U<�P��x@K�|}�u�dbgy�2�@�z��{��rE�1\S[/3m�%dT����qT*�1�y�Rk��N��QkTt�ӟ��yR[�x���������#u4:��\��1&?��2[*:=�'���O�!H+�7�i���V�e*��Ϩ���VS��x�o���D���^�_E��m����'O��EC�ǽ��<��]�Lh��{7��N�,EC�����N-R�V���!Y���DiuM�nj���Ry2��<�iP�@���-t��#����'�m�@Vo襧�V�]
h���<����5+�ϫv�'`91@Zx@o㷱��L�j�S�m'K׏>+FȜT���b�>]k!">̹~A���Aʿ��mZ��f<��y:��bDb&ՏB�c����E��C�&���:��嚟��v�)ġ����hy��-�e��J�T(DA ��f�x��J8������o��c��T3���]�=�]}.�8s~J��Mu��>(:C��2y�<7M�P����9��!m(�M�Q'|B���j����`	�=�����G�j2Ĳ�j�S���-F@������w��$��q���[u��x��R�U��Oj�����鋨Q�m:�N(tr� �w�z�����f좬E�D]�+�;�1V֬Y�f8������5T�S�̛��Q�"�vyg�Z�]������r��DϷN�3������b2�J8��W���duvY�o<��-�F�Ƀ7w+Qc��.��4pB��wZt:��YA�|~��*�Px�*�/s�W�������0$L~/O�X�PM�.�/�Ȯo��$��-�HxK��g��k�Kp,2��=�Ӣ����T�N�����/`ŽMv��q/�f�tȑ�(�F�a=5"�lR˦s7��Op�pQ��u瞧ݮBX����t}"=vu����Z�o�� ��#��	 O�W��Z��?3����Z9�z��i'JV��}%i] _�@5r��F#�����L�"ȩ�Ͼ59��^-4�@@�����q��e����-�ޏ�23[��|O�%r�^K����ɝB�j[?!����1�vE��<�9���Ȯ����y��t�.Ü����ip}{��}��yf�H+����eq���6�f��_t#��VtжE�@G�*��E��9^NM�14�a�tD�&���s��8�B'�i� ��q�s/ʔL��2��p$2�����[s���5�؂�A}bw�ʜ&�eFY���*���I��"�'mso�>h~`���a��r��Q�!��ܮ+6��T6�1x�eݯ]Ŕ���ti�F�]�zp���L��H��'ܘ4��7�����e�F�g\,�{�8���5�����d���J���~d�-�W&�3�
$h'���33qԻD�cu�@�{3lvt�?��]ؐ�M]�%����{{G�?��(2Zr9�i���[���n�o�-�_l����0C!Ў�(@������96C{�g��ɱ�%{�7�3A:
�Y����L�r����uR����d���+�I3ڥ���HBBB�7O;l��d)N}y�� �{',x��D�)� �)�Ϋ��!���d�=߼z�[���>iL����J�����p�F'u0�u=����/��*W�<*��#A����N=5
0���F�p�P.s�#���jt ��V7\�2�2k��
��. ���E�SVǆ�Ói=�4]��ʂoGH7���!z�݊��~x5� ��c/8>�_A�<���|���v���D}��e.Vd����6��ܘ��t�1�w)m�t�v�Dt�)��M	�&/H�M���t�G��+�_[z�<������
=G�Z���_�w(rgA�Xԙ��;U���L��m���i�Xoc)��l+I���~K��O:��'���L�y�S��\)�hZ����T���i4,�y�YQ�����%O��%�4�����x*��m�R��!�A�����ve���Э���"��N�!����S%���ۗ;�;v
z�=�5�h���u�
���� �,�T]|�&���䟍�"��~E+}���u���Ag6ZO\具h�x��i�y�8�fV���w�3�8�1�:�u/s�&xç���,)�=��B��)f%����	8�3����=gU���
�����BNL���ӧ�QL ڴ��t��zέ���E1�K�1�')0�ъ}�MC��q���r��}[�,l�'�>B:�2����ay�0�빌��y���f�`�|��-G�R��lïX*��Ԓ��W���/�����H�Y��3ϱ���vm,Lª�k�Y��� ,Ue#>}(l����l�˔��s�N��e�O󈀸�b"�o�H��.L�-o��bc�[�N��ʊ����\	jh& к�Q@�Ъx��=8{L�����T������w�t�8U��.�m�g1�3���=Pֽ��V!��N ���I�T-���G�A׳��H�Ik����D��fM�]� �ʍg�t���6�h�g���tM��X�]�)�Wz>4]4S����� {����fC�%����=�� L���ӫ��qMIt4"��U�x�7d��(�M��Ή]Z�:{�l |)��I�` e��n�����c�������Pˋ�:��ˉ\p�&�h��}��5�!���*F����Ĭ��.,?K��ƾ��I�ߝD��t4QP O���7�=l�Cy�g�=%�
�;��ɋ��V?�����]�h�:ݭ����	�'���dzY�,�8^G{HK�{xM� ��;�a�s>�1��t5Jy0/h�<J�d{t.-�l�����:X�W'/T��tqn������bUR���J�E�盜A�����y"�M�֋ܑ�a{&(}�X�z �Ҍ����l?�*_��ڂ&c���
�˸��Ǚ�X��H���j���JV��Té��6<L�ci��ρ���3��0Izd��:7s�N����v?H�?&F���}��ȓV���R�����N�bL�vp�� �����m�Y-H�O'����h�2�gDI���w�O7x��/f�򤈏2=3AY}��ShJl7F�f���/Q�t�l�)� �99/G��Ԗtֽ�mjI��:�?D�QԬ�(�b7�������w�'v��A(,��R�9����'�Q�j5���ʩ�("�_���LSP��o1�C�_���鷷��;����E!M)mN����"E|�Z7%W:��V��C˃�0�����ݛ���iG�.���<�O�Z��p9��lf˽��b�q<;�n���i��7�����7<A�����ZFf]!��"�������h.�X���a����0j�df!ᒼ�����Y�������k�-w����9?�y��F�deϖ���|iGq9����N)&gX+-���l?p��I����c���H�+����E"����m[nE�=BUaM7e���t�(zghu=ǒ��7�r[�$�o����Bԟ�*�#ZY�ڜ��#���]k\�� ���qh�  <Re��07�F*�_6�h͟�=ĥ=��%�*(��ź�P���s�y�]�!�sCu���-�����/��k7k���O��s-Sw��z?��\�������u���MK{�M��d��A"Y`zמ-uA�0�����.PΖX@L-o�a?��A�1?-��W�z��&�{������ �v�R��mH5P��`"VL09ɯ!��n\ ��B�������i�'Xp|`o��d������S�'s��v��l���C?昛hR�� F awP��k����`'x���:bRs�߁H	����6��Q)�ӳ��/�j���l���Y}�n3�w���`Ht��I�#���}�_��-dD�8#�h�9,ݭ�$��<��P�^���5L�/w�-U�<8�BK�)�cI{��09���=Z�`qKߛ\�0j���h��X&Z��L���0��O9���(Y[;,�9� O�C?6n�29_�������O�!�UW;���t�b��V',B'�ߴl���o��V|1)�{f�\�^ Yp�9�}���F��h�p����ؐw�������q�nGe�P�􇲀��S�؆ �חSǽwm�P呤h�"���\^�c����ݰ�/p�VU��2s�i##�٣y�xa*�˚�E&����g #-��IW���n��b.��.j���Bg�	'�n�#vz;Q2�<tE�EJ�����e��K��Zʪm�1r(��g3w��1=����	�������2<M9�Ē5B�)Ӊ�� a���L�O���}�p=�*��9��dP!jzt-�KL8�����q��n4H<�[���+��?c5�Z��������X��^Ɋ�(L�Y��"�S���0D���V��O��KsR�tH�°�Z��0�#���ƴ
g;�yw�X`�ĆL���؜&���e�@�i�G*�Ǐ�}��`�9��z@}j$�(�x+U?]�t�Z��q�^m���"`��o ���0��m�l��@�m������&1�(�9/Z���*"��O�TCPk��)>R!¡�Ga�U�^��ݰ��M3�Z��P�Z$�pV�JlɌ Wh�a�ZSe�l�U���s$�\���B����v
�^����a�����h�ǡ�&C�(ꁻ'r�{�Ove�>R�4y�T������."����q�%���p����H���օ��I���I�?�1:БP�׊����~>ȉ��J,_+�.�*��U�����l^�_W��@��I.X
2M����ǂEnq��y�6�.Tz��cG߬�B���$)��� @��#`gfF\2Lq$6��0W���F{�iۺ�']֮3��h��}� ��-�ϐ���灔7`��V�1`����w;:���3�!@y�DV	�Oڲ��w�$��<%v���8�:��󖹁L`���c�<��m��N���t���ŹT\��}V�
v£(M\�t

�rx�e��H`��F�y�:�'�΄N�4���q�����?����f��������څ��b(H���|%�16�z�y��E��'tS��]���%G7g�_�W���!e	�AF'&��W頰���	�!?oq�"��8�:+v)��/��M�ζ&O��^�4ʖe�Z������_���M׷�$����Kt�p7L��q�n�X�z�7��Vvp���x�m1ୡ0����AD�$HRo:n*�ftG�fν�\_������j͙q�E������/c�_��E��E(Wt�������ؽ����o�ꞤF������W>�� N���4�2�����%5�����d����hf|B�,.*l�`Ӫ��?�{�/�KA��&��輹�N{��i*Uќ�	��׵�o�� �Y�~�v;�hĘ{]V�~�@�1Фj���5��4Bx; �QX)��!�-�vɘ9նAv�\��C� ���Fzi�R�F�b���pǧ+;r�t�D�ՙk�''ZyZ��Jt5���h��nT���Ŝ�ګ��Sb�ֿ������-�-�OQʧ�$1���!��]V����Y�L&Z� ��j���;���|��n�eZ_���y��A�Q�0�*2�8����c��*�F�	JP�<^�
�OQ)���s�8���&,��L�P����<�����(�k�q1��&�z���u7Hx��B�X�+V��u}>��$7s��[j�	ƲE��؝�I)7�rp��z���>N͇W<��l��SV���ci͈J�[݈$B�B�U�mo���K�L�Y�ϖn��5��� ��6��T�*��.��2�:�'˽;�]��I5I�/t�LE�AO���mi�S'��Y�o
}*���������ݱ���'V�BO�Zg@�\
!��(�P�ĵ��+fm-�t�sw����C���Y�	�r�D��մr��R�B���-�q�[�j�Q���Xy�u����D�˃P-���?+�]U�6\0��-�&n�q%�϶�hНFv���O嶚��1��\�`�[�ReT']9GG0�����-Q�}�r�!��F$|�/$��=��D�?����H� ��;闎���i�����>��7{�7A�N����j�}�*Ӳ�zJv���@bmuS�~>3�y��	ܯky׿2Ģ*�[l��M�����O��|,��o�X���R��$"��e�)�P�L*K�����4_9��6�~Ղ�h*�����S���
��������:Y*B��L���ͧ>��������+��"��QX�d��aJe[z&��L��/��u�)x� LԓX��ͳ[ga��u�@�T���f�13��Cm}��7�!I%ݾ����\V�n���C���Ʒ'ȵ�˭=3/B&��%ː�N�����G�_�J�gE���_���V|ŵU`ό.�;����Fs�H㡠��i���� �ee��^�B�测d�B��1f1���T�S'l�.���]@��T����  㒐�;8�XUTq���&���5��vyp Z� �Ԕ�_��e�,X Z?�l���cH/�����S��^ր�ˍ��"����#(ks���m� ,����->���[��j�e{�%~��"Q��>>C�Am����F�&.��Eǧ�x��L�ep1�q80g>��+>����UH�����"����Z)��`F1�	��>2&w ���u0�@��4�F�S�Ml��уj�1:��P��F"���M�� '�^��F!����O�\��T�v[�q�����!t9\c�-�_�������is��t�Y����c��U%��d.��3s�����kz�����_T�QO C��!t��Yw��i$�B���8�;c�@�;���hef����e��� [eEq���M�*��;�U���`��}Ew������ɡA�`����ܮe���2cX
_x��班h�C�ݣ1υ��~#�Ahb��j ��7	R���ޙ��Q+d--���U��FFǋm��:J�)���C`��yGZO�(�0�g���@�ҫ����>���pb׍;���_+�2���z���bA�D�%�,cE��9��[�(T�,�h��p!exA�gA{ z��?��8����J�S�7�mCv��,��lS%�}6����8�=��5^�U9L �"+I�5��Ac�d�Y�S�wC݈ķ�C�j�c�2�	� �j���$FB��Q\�{���a��՚	y'1o��jx�Kv�NϪE�ץs��Z���.�������\�B�k��6��'� ��m���ϧ������'�)Q�Ժ�6L	�m�6�c��f�f���Ro�A�&�?���D+>wr��P�h�SHE��^��Q�Q�
2��6��^Z2bt�W�k�%T��bY�d,��&�f��_(r�kd�a�N�d����Y��I�3�M�$Q�Y�NN�$(?:����u������:�D��!8;S�N��^®��]j�;�_� .�pT.�P�r0�v�U� �h����6h\�NC���&9�����1D�窫�����9
a��zg�p����ɦ�����V^��&v�aSO��h]�W~�������8���d�Wn#�׹�����e>0�����wd�k��Ι��%�v�Lx 
��΀��R��&�@�4�o<�N�b�N��+Uk��hL������5���!)(��v7����;�5}�e��)-���L�Lh��K@�%���=sM�D�W�<�� �2Z��<]�&aK��!6L�c���
	)���i��ˌ���`�7�`�L�:l��J���v�P_ɥt��C�JC�<�b���dj��~=<��Z�gՐ%�Hn0�Hkӥ���q�\�N>5��>-���?�K�+�$8��Թ�^�6���M9g�Y ��G�F?�C�R�4k�
<P7'�>$~HI=��$���'wӼ)D��V��|$W#/�d(cKE��T$��c����~*Σh��Yw҆�v�V��H4P_�3�Nm��ll��&�_��aq;<�g��5� �X���=����r�ޘF#0⥹�����
��[��@''B��b(zD�s*i0\�Łx�{�F��k5�<��X�A䟛��Q�M����caE��Xw*f$���˙�3�|���OtP8�z�0���ߡ�5i�V�G"�qk��(� ���6�G�R�F��{�o�	^�[(i��wI��J��O��ڿ��2�ݣ��`��4�.��t��
�l��o��9��~�z�$���Y]�8Uj9#5�����������gM��6F��8+��8���Q��Lw��U]��p}%��Ց}�,*?�jvX5���/Lbփ
Y@,9���`^��-��Ϫ�ZܥD�;.�:G��Wre�B�7�������Χ��1$%D�=�	���A8��od��B��aP_8S	I<$u 1UU����bR@r�F7:^����ܛ=f��v�����T���_y���r��:��g�H_V�xig�<6��Z�｡��̣���n�I�����n��	Jʾ/�=i��}�}~��3�n>T�8k������5�k �5pЩ�����_��`:�(����4dR�3�p��ؙ���P�^!'��&� Q��cƼR1����T�)��}�`$�����)���q����'�.P��yu���-���h_�`�&A�����s����5�~da5�KK��'n�_0N�}�����|�9�l���r(�k�׮�!�ٿi�ye���ј���}
�"N.-QN�t3'J�O.ļ'��qe�~���|s�Yc�ԗl�7�^�p��ٹ��磺X�G��6\��"*��Zw���蹐�!��6Ւ�~o�ys��Jbu�e�v�y�U}������_~M�����+hֲ��Z&���Z�ODU��m�	�����s�����ƙC����$=�:�WѾ�1�3l��%[�Ke�fz��S�ڵ�oCuN�r?{m�I`u�c��oĆpڐ���ƅ�����Gq+n��!�L��-D*6=��{�1�g�XW�6��RI���|�4�A�_H�4L��i�ZˋX���@YV��Ɉ>�}R����*�Zh�}��uIr�C��i�����	�;ǩ�GEy�[<b�RT��׾Y���1=�K�8= �wQ�B��L��;�7_\l~?�#����w��?��j0�����{JG�� �Z�;��G����4�S
��L�ّ�&����m
�߸bT��}�?�=G>��5�5�@f���U�\u���c�w_:����OI�/�k0���@�<V�jR3B�ecĕ���]��v��b0וX�]�D5m�*��/1���	���|��ԃ\f���8��r@����U���+��%�qO����ǖQ�(ґ��[�'�[J�.�ΓC��˅T���e�SAS?d"�;����#�8����/"��V��a%%YS���R.iI�D�P��c��M�9�*I{��T���6��? l��oUo�H��F<������;!�H�HN�ᝄ)mł����$	��?_�R����C0r�&/�
��0���RuB{w�֍ce��R�_4��W=��ؤ���w�7�7��1��Z1�/h�x�P�S��
��RM��:�f�;�h���w3zBU���WQ�j[�	��G"�?���y8�������X��Mv�Z��v�1�����5�3��y���g��L,�Z�+�B�i���UWH�<��:f��Q�K�������]=Hp���޿[�ߓ)�?�=�����1s���x��f��o�I|	���kZ֎��bn8^}��a#^q�SCD�E
�$���q�xKW\����~rv~��2�Pr��O������T�p�>ry�9G���x}o_�^�So��A��Mm��\7a@�s�4�-U�:�ƩG[���-p��n����Ҝ�}��`�XM�>_Oj;�ؑ�O�t���K��^��TEE}��wc�$��L�D��P�Bߣ��L��P��=��}G��p�At��&\��d�Y B^��l���<��������`�r���A���_��0"~��6"��k3�]Ηg�p�-��g~ݱX�t�I�"ѻ�1�y��a��@	��6G���
+[ْ�-�	�<C����v'�����n��SS����Ig!�m�d3�b���%��8�<�/A;[��b��,Y��tȅ�/Ů���N�_�^�-�4�rQ�V>Q���K��Aoz0tE�<�d��ַ���(�O#�>� ��t
ς�j��VŻ�Xd�� �o��n���>� B��vi6uM�����kB��1�Uw��O��sn�P�C�E�]��-��x�g��\�E�]2J|�B_�5�~>`�\%�Ν/�" UM����݄U�ː3�wx�dl�oK�ơef	6f��8k���6����E'���4�
���aˎ�>Di�V�
��XM��Z��X����ۛ,��t������ď�UO�,���<?O�}�(<>��,�4]^�v��c�lb"��t�*��r�b��C�������W�(W�y����Ҭ�%���
25��oGB~�e�Tos=�hK�%���,Lo  �,��O粒k��k<��c���?Sm���]�������ي�%�̘w�p�2�߆�T*��
�F��β_iӎe�����~��|KG�B�@ N;�e�~�=06�2i(�Ϊ�?� ������������$��o��+������p��k���Y2�eC�:-; p�;^Y �)k�Zl4�P�(5��!�qi�� �D�Pi%;��m�}
&��������{l�g�v������?<��*��'� �A�,{�-�͞Jq�����^�j<
y�s���j�<
+����Y1+&t��̼jֱ�$'��]��/I�@�����&A1YH����>�N��m)r��B�!�����{�]ջؑg^����
��d+��*1+�~�d�[H�h�<�����,�j���@��O�w�h#�����;\�ޅ����R}�%��F9�!3��.��<�g= �	��ߎ ���w�x�:^�`f���'�B����G�^̽��!��V�/ܪNe��>�m[��W�{W�Ycxv?T|Aʵ��kL,|��[)Y�L��#�����ì��q���w��� ����>;��
q���[��ʁ��)T_p07�DR��L��eJ���=E�����m6!��"ce��%a����X�/ζ��I�o~h�SK�`S	���`5=�|�JgP���T���S?ץ��6����#{���Vk֙�w6���8 j(������Ȉ�j&��4츠��	������M����f�����ac�o�@��-�>�􊇑�Qy��@�[��g�	���m���ᰅq�Σ�f�¿7J=׎�����U-A_,����������n�PY�ώ�ԣ���ڜr1�M�-z�LY�;�ʂ��Z����1��F��ZT��"�O�W���E?悜Y��TZE�I�W�C/ݫ��^0W_��o�3�;2�U��[q�O���nPT��R�Ҟ��ߓ[�S�� �N9�m\�8�l�?�+ii�߹Z�9o���cd%�5'RJt�V� hT�E��'֐(�y���!�C�~>?jIW�>o}�� �0&e��r���%��Z�=G��z���ی���8&?��r� x�F��C��k���D�c�?J5�ӏ�'.�Nm隑|�h��Ǹ0u�����{��S�,X=��Ȉy�rw3��T��&D�0�h��}@m��˵��Mˬ���<ܰ���qz�V���b#۾\��{�^�8��G���<E]�;uٌ�zd�a<�����f�}�u���D�(կ�ӈ���W/���zX��:8|n�?��Bw�~n�+��s_�ib�s�O�S09�����%M��ب����֊F����t�B5~̀���~�׶*�`o'

��v!�:;wb���@M<xi��3�K��i����d�tJ����2�hi�,���\���`�_&�m�����z�8�VT}/Z�����[�-vMK��%��)��� ~F�U-�?����vK��ʛ� �emG���V)0�GV!��ߎlr">�4�O�k�w$V|wf.x��[����X�l�[8;���b��/۶2��E�;8��j�H<S6�l��Z��	$	O����9/�i����q{u��`n���$�I�ӂ�YMv�a�jHbhƧ�֫�ke�b��Q7co�~��h��rP#�z_.&�h9kU����q������hƔ[�h�3���r�r�����Q�Vi�ok�DV�,3�|�:K����^Ёpk�7�wy����N=I@��$@'o��I�1�P/-K�>
��+׏4�iQ��aA�÷���o�=�S�n�a�ע'�����ϥ6���$n*����c~�d���a�8��WF�M��,Sȿ�'!�R�FϿ�bm����e�O)�]�f2�l���F稽T���bt���j��F6[��̗>���$JLz��HPdL��ǿ�p�Ty�o	��|s'K$�� �(�5��e*$�/��N*?�X)�;{0�r��6fw�Z��ea(;����~��ԹV�f��9:������Nt��၇Mu_q$ˈ3��l#2���2��2 Lz�)U /;9�d�g�p��DM���YU�f2MF5���9�h�M$����$>#�H)q~�t��X�rɇ�ct��r��P4��BD��&1|����T�c�f����܃�������X�\������X~Ch�"��ъ�'�j��D?���Մ��92^�~S����B\3�	�J��E!�����3�+�%���	}�w�@���W�RV��5��z����4�,`ٞ���:h_�a�*6uo����Z���uX	�^V�3��i̠�?�Q(�����?�m����t��~���=��b���uvTh�30��H9�㮿Aw�6�_�q2֛������NR�0��'��F]������&jF&ȫ81xȼ+P�	��O�
w������A�����;*�ۑ
�x)��ђ�� r��z�\��"�ff��r�ـY&�Չ��p[��hǾ�!�'y:D{�ő�<����h%lSA졕[��+NW)E�z��B!�2������_�.bj�較8�ԧN�1P��;��E��Wɳ���!3K���+z��y"�ڌy� �k
�Oeg�C���W;$�f�ˤ�Ж"��4���� ]�Zr=���Y),�sjڤ�+Ĝ��5;���N�R8���Ie�i�������������g�܏��rJ������S3���ܗ3�K�n�%Ln�t?����ZT�dHŷtnjG��T�W���*a�:̵�/��4>L�L��{&�a�]L~�U�D�~@L�l�,��[ �LD?�s�uY|�?<��I=a�^�4鈲�E��Hȕ�T0r!��c���%�6�q�&N�;��B���,��=P���	XB�K��}�����d:����g�mx�@}�_�ǲ�q��B�s3�Gλ ��+�=<���&�@�A�m�~�8]���X.,g�g`<�2'��\$��5����*�<�d�7$��C��ي���"�5����m[Rn����ϸ�����J���v�����ب�BZ�Y��BQ��"r��#�^���c�t]��8���u%+,�wy�k����FTCtۿ��&C_y�_k�#�-��)������YRA5�D�z��M*�b�17��1@�p�DZ�o4�4?/��kي�����}���J3�[q�o5����o���#���c_���������)����|�S�)w8��=�F+�GZ[$u����aCۚ�f?C=ُ٭>M�hoڹޠ�K�$1[��};��!-C��F�~
�8D=Q���[����N0���絶��X�32����Z.1��x��A�0��'��I��
nO��Ԧ.�8[)_��@�U�k?�k�4T��9���'�×�;
p��������	?�/}�ǝ!�d:�wr���}�EP]��cUW4��>�t�T�|���$h����R�5jYf�Ch`E"�d�!C�}t�(�6�J��p�U�[�%�������A�'��̮+�;m-�cQ�EW=z��4�޻v�|cþ�}x�aJn�5��J.��=f(ی�LT��p�����<�䤀�S�}���))pڔt]�ʟB9'��V^L�6���ꯥm�˴�	t��q���z��,-?��C�躛��,2��5O[�;�b�_$��c[;��z����	��\�S�%Z�6Re�}���� L�]1s">#�Z:�#G�L|I�+�?��g v���l�������Iޚ歧���ړ5��F��n�*!�j�)��"����p������l�"f(m�n)0�t=�v]a_���mU!�F@�q3NsZ��E�SIj��E	P]�LU��ª�O����oz��,~�����
�L�6��ZG,|�*ԥ�/p���kv�Q�*����F\B{	.B|�=.�"LE��)5R�e�.�|O0���=k��.����؊j�:�zD��C�B/�_�=�
��~�h�),������iҝ`���0hV�i��Y�Q6��T�n�;��_H�/��4M8�O��/~��C��n�_8���{Wl�H[13��T_�Z@0TkF97��Oׁ�����V�b���gg��2	W� N%��Z���C��%�yN�纟כM��Z#���d�hQO�n>�&�aDT�]�N75Β) Ρ�&�m�z��*���s	���$Ц%G �n�=F�r�"Cl�����Э��0#klc�X��J.�cn��������X!]�]ɧ�2o��yG�L�t�q'냯�e� %��W��Y�x ��3�8X�#�O�o�$����)�CJ�K���FY[�{Hܯ>*[�o�;vrNlE�wxlJ?	�!%�$��ޤ+Fծ�Iۄ��O
[_>�cYG^Q}�Ϻh����8%��j��MU3��7�g��/{ �*���p�j��!��8ӏ��H[+ZZi�؎�%!��!�($�V!T�<%AK���0��IY�w�$�e*�]#���]{�w��YA;]$�}f�m���7&�ea(��^>����ʅ�7�9�lj[��~l�"���=ȩՂgN����3᭎I���_w:��$�i�`S�������3v���˂5�0�t/�(����Pf�"o����b�rt4�%3m�F�9�}��P�t.l�������h'6$�s�z����.~�4����wqY����<�z�;h��~"[C+��<�i�ӣ	����D� ��˱�ڲ�v���`��U)������V#9��T��؁��P�;߶��@�W^��4�=���Q9����
/uWLm���h&<m���C�8E[YK���o����a�h;�RBԵ{}��b �ۺ����a�f�݂�cЮ+��@7�'����3�!�ؑ*&�$0u���;''I�-�Bj4Dk5*�"�O:=q m��������ޅ��.�7��^�f���t����A�9�/��@#�s�]/��@��,��/��v^���3U�3s��'G�-�X??������\�
߃�=�iqť�*�`��rW��zs�����m� �?��x2{g���#$�z��ڧ�"�C��nc�|`��Yh�n(�'����V��7���6&�:��7����'�m�7��O+�]�G��@�m��V�+M�@# B��	�Y�ht[@���1_C[A�TĬJp$������8�8m��Y��\����j)�9rp�5_�	�Aod*�YDj!^���ZN߫E�q�t�ٕ��@��gg�0PRM`��>������8��g����DfM��:�r�M*�p���f��]@�N>���Nא�B.j��)�M���s<a� ���jMb��b1+u'TGd�}s��G�PQ2�&Se��2I�[.�r/ߛ�8����f�Oh����x���|���4�8Q'�Zl�C������M�8� n���[�۱����
#Pa�T	�ҩ�L��N������&c��&��e��S��a(�	878O�����N���?�.��U�%�2�������<�'a@@�C�i{S5hEu�"[z E��������`h=�����9��ZIs�r`�Z�j\��k�!�VoV��-���
�V�����3����V��@E��G@ꛅ$.Wq���Ys1�ok�[�	�l�e��I�Co÷�Ni��%��j�x��s��;�١M�k$�5�qNm^E�As
ؕM[�h�fMD������D/2ohԪ��:\�B�%8D�FWo����p�F�M5Ώ��ӏ?*�T����M����t����dO���w��2���%軠���݋!�I�o�^.��Z�W��,4(��	�"�������B���k6G9t^�5��T��GU��3�*���t'��O�*NaI6���Y��w����ͰO���<��'�%N=X;]_@��O+�JW
�=
�X,��0Dǁ�v�A�Do�ݬ!�z�:�48��`�6̹m.�$2!#�t�f��*��ۈ�ã�?�yg���1���m�d���R�M�,��-�T��	 Ӽ�5,<�)�k�I2I�٩��q��G��+��4ku�J��Q`E��!!���E3�B����G���C�<e����_�!{*���Bf9eG�h�չL��Xd��`�d�=����Ю���)u2s�OAvXE�Ρc�?Eo0)�������ZnJ	yl4�`����f���l�N���W۶T(�q�R�(��u�����hn�������y�3{;VzO��%y��0J�Y�=>ʠz�T��������	ØZ�Q|E	�K#Yy��M�u�{�C�������?Ǐq�B�Q�x�.�r�;\���]�AMsmS��zO����ɼ�D��K�!�\Ѣ�Qs_?��π��������+�n�_
�	�a�8O`v+9���(������{��HXKr��DK��3�m�3��׮�%�B��$ԗWv.b�����yjHjY�(��d� ������T�)���ɾ��|�<^Q��6��s_~��dT� {�U#+Q�lו��\�
�|�-.�t:��}]#��ď��e�kK�řj���טѳ5&&�h��)��5r��PC&�&�Џb��j�jn��{_j@�U��D�`�goEt�Zf32
L����� �c�*�rlco=7��1;��Ꮿ�K� eO���Q�D��Y���Puf�<�x�����-I]@��[3m�~�����f�!�	=��E�*��e�H�{0r�����K?
�5��S�*�����-4>��p�:���?mͳ)�'|H�ҥ�M*����k�p��"��_N���Fb��m�>l6�.�,�Y�p�0�A�b��/��lh�[+3�T��K�Z��L���i��̏x�d��A���͌7�Q�!�PS�asD�y[�MA$aT+/M���C$�dD�v��R�F�b)�n#������ƭ:�ј��塩���5�5�uI�ڙ���*!z� @�Sm�9������y#���$L��GjzaԂ#��:t��$uE�N�u�%����A��r��ä˫67@9�\��k��m�tH���Ƅ�W��3=��#�۔@�jh�?st�1:���QuNΪ=mD�1���/���M�=�G9� �:�L��	.#>��:�����	�8[����V9 ]HN��_�gz�s.Uo;����30f��ݹrW�$~|�W���q��t�n|�G/��&iT!�Ď/K���H�~���<T\Z��������5�/YQKn�h(K������)m�TR��� �jY�C�v��ڌ?ϻ���IJ��R�w�&.���&p+/�����ե��?;(|ڗr���W/t,��[�[�Y��PY�ͮy�^m�G�+B���f�%�K�~�qUAwܘ�~�I�z`r�[_}L��~	��W�r�6Щ����ꌧ��hb�"�Z��]L�@qX�)M�bC_zV]TD�F��:����i%��"�=������ÛV~>a��ߌeF��)O�V&
��m�L|
[����{{��(��.��W����+���@�����ߏ���U�M(�Q��ڔ"��${���6�4�#�lCK���R&�As�~���Nc��2��u�N8�.�DB�v�^iW����饦���s�~Q��=w��%�ǌ�/�*N~��L0���n�
����"����>�%��V�qe
ۡ���K�2��.Q��� ��3��8bY��r^z�7��=Z�:n8D��st�<:�d2��s�ld�8I��g����Z��������[8���Ϝ�~�X�$�k0~|ymP�]{;�*s�K�ٟ��'-IKs耷�ۃ����0W��	P�)�X�s�u�m�r��B�'���K�Ql�Tdx���qL�a�ԑ��jh ��"aHg��%���k�nF����('��|����qK~CW]�7����k7X�Z8�?!����y2�n(�"�2w����-S#
cx��)h��t������'=u]�؈Qw���<e�]9�#����[la��G�P���.H�AO&�_���h�C�X<��^,ڃ>�׉�;�.P!�w	�T�j8�{6�G��ͥӀk��7W2v��9+��O=�%1��{o�1�ޭUB��w<�N"g�U���R���
ʡ�� ��:k�ǟ�Cd��i&�g��c�[�"��I�ŇÉ����Sx�_���Y�U?�4�����	�\�ACAL�P�w���7#�h'z����ԔI���AM5bj�[ ����� �7���z�/�8�4>������)BiH�J����5�ALBEt�Cs��鄘*��.C8X���a�C��,8~H0J�NУd�{Br��ݸ5��ru�����*��%7
�´��c@��<k�3/�|�=���9;�$�U*ßg����P��GKM]]BgRШ�K���D^�Q~�0K �U�V��NHTƐ��/ :�hQ0��i�D�^��A�wn�1���ў{6!d���u����K����YZͦ]T[��}������Kg��r;B_{ϩ����j	3���Ό�T](0���T�EV��!.0U+�h>���W�Sf߳�T�b\��-�����*��3w�tXl�&�rd���xaǍ�_e�����o��Pi�rĠ�r0��<�`@ �wj]E@f:�V\J%�%��3_9s��D�&��,]�,��Ժ�W�ָ6���X�+�'l�~�'a5���/e��i�̖$�7	F(*z��J��7�=�R�[�G9�,@	�bPO��B�qO���qچi*_�d0Z~W�}�5����~%�B�v6��
�_�����K~��&���Χd	4�����Q��+��[�x��e0f;�'n�Uz��iM������M~��u���2&����k�;�W�9'Q��)�����5@�[�4jPw޻��6�!���%�םr���r�q���Z3pp�Ni�u��F������-��9�t�mj�M��+��2XBz����{P�P��7� p�&��}�� �4w&RX{��46"}'��Cb��79��"�I�?�.�.(������)/AE��qjp��$Ӳyq�`���D곐���`$�Eݑ�r�j@���7����9�ϻ�o's���5�n�x�8��Ue���	��-�����ɩT���g�N(�i\���H��Nz/hSNJ� ���`t�7P��C֥�/��&�H����?t��If�u#�Sp�Kb�lI�s�}��.e�`q*��?�?WyroB�U k��<�%0	�{���+�X���v�y-CWRT�YRj��WI� �ko#G����yKU�!ANKSԒX;��:l��'C��jQ�d"�����
�;�1��} 5�D�ʍ&5優kƘ(�Ql���z����O�Q���u���_�	*�׮�%^d�-1h�b�0,b�T�2�tӛ�,�|/�E�m�qG�U��̑�	�}TF�e4"��m�lЏ8�z	��D>4t��I]i�-b�]���LV0�?Fs�_N97t��qPi�6���@[;�͡����ۉ@uUT9@����h�˿C�UBF���w��gKh����q�8P.xL��B�+a����>v��?��C�� W��8j�Bz�㳢h�ύ׊:�(�=.��� o|PF�Q�=PJC���.n�R�!B�z|.%�g�@�D���$�{�[(�r���ܓ`	4�FH���S!11�FZr.�3j`�2��]��&�M��1�����0Ѡ�7B�ص/v'8*����7�*2��8v.�#8���NB��wxu0��r̖���գa���,�\�VD,��$#o櫔EߛE�]���ݙN���4ϕ"�Rf≁�7���?^�{���I��4�sB�Y��{�E�ު����uE5#41R��>��00oB��Qڍ� vK��G\l$W�F:b)�k<l�m>/JJ����jJ���,?ۺ` ��7���~�\a������>m�bA~7i��'�m���)�"U}���g�~#ew|�D������柿�!D���QP�
ȉμG!�Ϗ���������W^��-c��3,��e�r�A�waem:�q��J��)����K�5�e��Za�T���"��N\��iE8P2lt��QT��Ε�PMx�=}>�ǭJG���BW:҃��OX)��by�dvk>U
I(�֙�OE)��ܺ�p9�^ȝ`�Q6d�E�<�t�[`���\�#)�rPA]c��A��v�:Ϫ�|5?W*���!j
�	���Ц%��]�v׍ �Gy�v+1���"�^�PD�}�ח�$�^"�D(U�h�ŧ&b�������<<-��%+c�(��2� Gb���ٿ~�9�/�&�?)���?��}����[�с4���P[e�.:��&��pqJ2���>ϞH���d�No��K�+��T�����piWO#�.����X�,QV�������9u6@/�?�>��EF�u��g�(��i�9qT���I\<l��Cղ�� `]�K�'���b�����_A�[��Ȩ��K׏��'�y�v�(ج�\y���H��0��ly��0�X}-��*�''
�P'8i*�fpH�t ����uPO�P�p�#f�wǛ���t�kV=��3#��:}��:X^_܆'���2�׾�
���*�����/<���z�E8x{�.�jވ��y�����Yƒ}@љ)���nA\��R'yUB�?��'�t�Ԧ���+H���|�Z����ڌ���0�:K�FI]����UcB/,�>1����(���T�Y��4C7�YA���"�Gh��|\fm��\	��ݳ�\���:f���fv*����/x�H���q	��tR)�:0��L��f��i"JEs��q������R��S����;���U�^t���.�-4t��.yw�F�Y�|���0�l�X�=h��D��1˩w�˶Y5�:�W4pĐDSpx>B3�Q�Y��v�� �' Q�.\p��L��`#5y���7+Qngt.(�7���i?v[z��S��[�
���"|�Q�iR��!W	K��l�Po~���6��5�=u{lZ![=��+4@=̶��2յ�!��|ķ��o�gq��`��?�"������F��y:^J��H��La�n��Nb�`���N`�u��n�?ͤ���b�¸���3�[+�\�ߓ7wo�#H^+�L������:��yI4Cއ����J�_7K��^��J��7�Z?l˾��Yϙ"#�6a���^[\��uMH�>� 5)޲_�o��#p!��]V��$��f�R�����,g:G.��'�=^�/�_:K����V�ჹ��-B2_�WVG���|�&�FT=�.���hu����$o�����+����Hxs�1�+�T,�%�F(��5T"������Ei���~d��d��ؒ�~��?�"w�t�v��m���1��9i�7R~J㇉Z+�˩F@��