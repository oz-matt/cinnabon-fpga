��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD�w�6��]���/k!Bu��s�B82��ɨ֎���u��yށ~O7u`����g�������Io�|=�K�\5�z��I��2�zm����8u��*����>$�?$��v��pw����C�r	���oly�5�M[_��%֔b���~��L ��Ƙ<�8��-<�R�2ԈW ����.����h�%j&��v
;�r��?] F)�r�_�8���|�,F��Lp ���d���q~������˼n��@x�&�,T���)�N-&�o �ߒ�@v��TɔH�PBdCO5/������L֌#d��O�[��X.�e��������I��;�����,}�!Zˊ��.�V�DN����N��
�� oD������n��(�v^�#m�ި-Il��*>tÊGڨ�DB7%��`��ϼ��>}����@�Z�DtⰢ �pZ���,��%+���@H��<��p�K�=��25�o�	��A�`�I�7�Â�Z�O���nn�w�P]�����п�z��J�!m!1�`FR��Xu@��������b�.�T���璚Ԭ�wd"�x7ͯ�-���A�;�^�	�I��41jI3�f4n���$�2oy�74����mQؕ!0�jZ�=6NEݮ��	��7@�Y�y���� �, (�BgN���������q�yyĉ,PaRy��S�5�)��^�w40Y_o���܍R�dٮXKb�0��}�P������t����m�:3���$���7�GA� �F�:�J����<uo���\(c���_�ܷ���g���ⱎe�i��6�-��$A�s#WbH��N��P�Ե,�ɹ�I>#fG��Ǣ���3��9�Z�
`���4���p���5_�7L�?�f��+ڊ%�J��h�n|N��hPm�Jf��M (\�ʌq��) �q�gD`+�s4��͜�'!G%��:V=+@3���(�l�U��>���P�z]dϯ�$�|�����i�RH��s�lRV�+V��>��kO��J#.�cf�s�l@��%q_b+z�ʛ
���,}��Q(�?����x�ͫ��e+�U�-Aa֩�y�R>J��J�<�P���+��՛�_e!un9w���J8�Q����4e+��m����b&k�����%=sǠ�@p�#)�^ت�����0>��bezv�i��L*������ױ
�\ҽ���N��>����9�$|/,騃��M�I���~ZP���ȥ(ȑN�,B�aD��Wsz�V�	�	:dß���e�D�����$��3��Mcū�Lw�:�Vm.�$]]�i�s�~b��	QK+X�*�V��g>�BA�N��}s���q9��ź#~�6A9������@���K��}������TwR� ��R$�v9ڨ~&O64M���]���95� �՜x=S�Z^����ZK>��0�S+ة<�\7!%��@D��{t�TO���gP4��m.Ə���	m����w�6�eWb���J�z �׊+��gϓ�`�Z�nC���s�T����{Y
Z�ԉ�+|l�$�9��H�x���O�訄���/v��#��X`z�S����B�J��8�#˷3��}b��Wm���#�����f�B�yY{�p��T�X���F-�:כ�h�����F$��0�����D��]dY�T�*�����Yز(	{tU*���4�$˯�{�Y��<���=�7��Or��H���Ϊ��[f2�O9&z>�1~{�(G��Ԯ
�C�u ?X0C����}���z��K���ʦ`���(�%|��ų�:����������]��>_�.���U\j̖?L;����E���x����\>P�hҢ��3Z����٬��JSMq��tDB�n��>�F���&R)W+�)��	��J+g��f�lq��PJ����sg^7󞳞5 ��!O-6�$�T�@\4"�I�$'7v%EydeC��u7����63OI<l]��.�0׊-�Kr���s~���죯T�}e�Q����#qL��kkA6���:�P��b��>t��.Q�g��T��Ě8���u?�rGiY^@���aFi"4�/ǌQς�w6Hг���ئ�����lc��)����2�����e��w�忡hƹ��G1�͏�� ���x��p]������̎$Si�6��&1|���f�x��;�H(���Q>�Nh\�y�c4�}�H�~�3�H.7ŀ�R�~��<�%쪒�M8���go.'�=y��F���RCx�-W�Scs�!b�X40��ȍ!��(I�pv�W.�~�(_���]��)X��q��Z!�}"=s�Q����r�"Q$\�S@��G�|欂3n����T�@�؅��l��()h���q�I�Q�+�تς|�˯�{�.֎jçi��*��8tݲ�H<b�+�P�g$�G��\%�a"���^�D�v�B~p8��f'���aQ�l0�|wY�ܱ���)�� =Q��\e��9�@9�,�'�V8��aN��%�����+8,Ō�d�1�ӆ9�cK�g�9��v�7�i�S5���=j�t������2͓���z�>Xc𓲀]'��o_��L]a8��d�&����C������B
��pQ�?��'�r-�as�%��q��o�������d����?n���>|JmJ�?R�	�K;K�+x���;�ͽv�+��?�2��*xI߅��?�6U!�۾���-�yXw���W��ԫ�s���q�,�^_amOm7�D@���^����)�n��H�Tv4RZyD_=�:��0q���eGGb�gю�扳�q���QA��l�# @��ca�kH@[S�܉�(��Գ�\�;��|�����i��W|$���p�7˗�Qf�S\BE�Z�2�PUs�FC�.թSX��腯����d�ϩ����u�]ML
���:S��s��������]�l{4�j`�:������d�7Q�SH�R����3��~�BVp3_ �<�gW�C��s�0;-�|�T&��A��2�Xql�����"�g9���y1>?`�c�-�u^����8.��h�S�\��aP�#m�B����[���i�Nq'��0�w)Ip,�|͇i�x�5`��}�k
}`��`�7>�T\d/	�q�T�K1,9� �N�V�B^�.�����9 �VV�u6�Z҈���ZRS q0��i�P�I�	 QhO�)!O���P%y�B���"�����9l%�`�]p�}u�H]QY��$��y��7��y��d�%/���Q��-���άB褄Vj��Ba"[S�gLɌ��jꝉC�]�A��񑗕K(x�%&@Җ�[(��D���%>�lA��8d�df��g<�_��!]55�&���L�
6yDq���<�2Q6�~����͵fޙ�/���S�'#Y���<���#�����r @��2G@��{,'ǯ�l�ů{�����|L����3&.T�vE2�{o��t%��6,����pc�Q�7��A�������3�]Z��H�と�g��}�R!R9Sޅo�r	�E��q@��#Y����ԋ��R���Xm��S�e�<���&5�3��U�Y�S�5�4�n$��� !s&p��u�X�+�]�Q3�3˝���HKn�7�I|�����K�"p2|�_�7�6D���D}��.�v���#�g��&5�O�+7c2QϨ:w�Y"y*��aw#[2�m���ϐe�����_�@���c�Gp��f+�����������^ѓԸ����%��v4��{6෠����:�7X�G؊/0�U8�f������ V_ބq����K5_5($��y֦���-�����\�&p��q�����hT�z#5j�h����"����?)�5\��Ǎ��t�:�wL���G�GO����X�ܷ����m�rȇ�$U�9Б1=e��Z�1�/���yf`��IY��������d�b��Fl8>��%�� �O�`hb���D�����00神͙͊�������#RϽ��g^�����VN����Ƞ4)o��~����ٖ�p��'t٬��9�f��Q�����IQۓ�<���}��X��!C�S=����,���s)�M��m=t/�h���fB/�V@W�䗉]�D?��o~�����&
ny0;�gm�3~���_Z�'����ߓϴw˶mi�ï���pj+6C��X}F��P�c 0�2Q�Lw�4O@���t�n��IA?}̼%"Մ
 ������2�nvC:z�\lM����o쀰4�I�Fq�؎/U���W���+[G�7��@�:��ۤ��>�p|핔���ߐ����"�|e+�&*y�μ�(�})5�G���s��ۻy��ݬg/w��W1���|�bdu2�"�3��E����?�n�|���qo�XȢ��5�K][6m�C�-����)�N��WQ��F�� �O�N��۱�a�����EaPqT��aTHo���u�?{k��������wզ��4^�N�Ƴ
*ކ�7c�@!mzX����{9��dL���R�"��u����'W~ϘSX�ϥ�C��b�O����r@� ъ��q
q�PXe^0=ob�ԗE{-��gT���9��桾���L)sQz���`h�^�BC���}3 �2���1T�'��e����kp��4�W{��8�Þ�ѿ���y�#����)�6�\��z,��鴇��5� �����,s����*=j����5�{�������c�%����U&�������8�6�0q��x�I!oQ�Z\6�eBR�$T�3d��p���F���"Ix�>�y����.�.�#j�.��0[{b�!Pg]�èv��DU������$�I�k�҄H{ɧmu� ��PD1���I�:
�۝�c�K]��D^���8�����#��:Z����%�WK���uG��n.�B���&q[J�������Fz+�Y��bY��V��:M,l��}y�eT�537/w��s6DM���ɕ��Eֿ�Z��j�� ���2�r7��j����$��U��C�[w�?�{\&H3XUI�)?��5r4R����+8�p�P��� �BO,rI�0l����a��J�Y)g<6f������P55Ұ2d�f�8���<|+��^����^�K��e!�\.��N�I����1�В�������H�2�f���:�0e�m��uE��#]<��o��0!�$ذ�˚�(��j~`�<ɍa�ɧF�e��3 ��Ht�~S+�M�5�+�Ⱥ$��OY��YIX� �۵Z�3\�	��-Y�`_��u+���A�;�5YK�s�Q��=(k�+�N�t�2�5�����k<T"Oq����59>ռ��,@{�v���`��`!�P_\�����$��k\a��w����<�+:X�q��ƻ���8#D0t	�1�J��+�l-���q�}��q�	yA3U��`���l4��d]��8J'� me��#Bw���Z����OY|Vq�o�8�>��S6Vƿ�[���w��d���W�⮉������4Z��&z�후��si1�h�����?K��Õ�ȹ��Q��K�-E�TH��˹�aK�y>^��ئ0�s�Y���ßʬ1�& n_����H]��Y��ʇ#�K>��rȶ�����.ɲ*C��9x��u�����,�ü$L?TƄa��O��U�3Ng�.nБ�]�ϹE��h����5m����>�T�AZ�U�����]=sVi���%���fSp�0�"�%4�N��h�Q(����4�h�ٯ����`�/�xe>a�<A���ݑ$�.,�T�:����͵���ٷ}�kVF>�/Z�ME�T�v���W���Ӌ��k_�j)3��G�&�;0��tm�t����,�-Y�O�`C�&� ���1��~m�4��J����h�HD[�H	C\'�Ne,v�r���N������r���PiK�;ܻ�r���1	�U*R��Џ�L�K_i��KM9δ��+�[*' ���q��>�P�k�g�l:�u<I6��ͤG�I5 =����ڨ�`Ag����&+�a_~׭z��]:��_�����5��<hQ<r.H9N�,l�&��R�n+G!��b��
�eD
:����E�g�F�M��`�*v-��!�����l��y�ԋ�Ͼ�$��\UZ�g����|j�Ƭ��翸*"V;�⢥#C�������J�D��pX\N�I�H��近So�.;��̳� ?޻~�p}�[r�
2/��II���_�Ωsmq�<Ԉ�(�º��6����i��Q:�5��!'!��_�����=�4��m����M� �
��"Wz�,<����uoV�彑9�͝����^
�Y�K�q�X��m�'�^��2x����.&T�#4���	36U�KM����}ę�2z�e�,�>�'�ᢽ�|\�iqo�A�W���Sw^��ɰ%/�=u�*߱��!�l�d�����۱�$�q���':�u����됴�#o=:ReC����&���C�]�����UI����X#V�.�(�(Q�/˭i͝p�c-ٯO�㘰{yX>N��/�8JZ��b��y�,�ۦ�8fp$:�2�Ul	��b�Kw��6�}J.D�_�����E�~Z��d7�n�L+�iC��5���劀��%ш��
(��l�݋V��q:��R�E���I�Ɍ��C;z����7]#�H��� �8�-U�{AQD���D�5<�('�
Vhs�@���'�C��C,ï�{��Wp�8��8a�o��p����L�TMD�r�[w�.������8q��������)Q�J���A�Ji����f
��
BN6ﲟk��܈U��15"R�Ѓ-߸6<�0*��9ׁRM3?�<�y�,�&���F@��T�X;��	���y��I� I��s壎Du����<��D�X���+k���V�g�8��o�ɲ
��w��T� �{h��,��jD�Բ<ڛO���측-vBf���x�;&J��ΛL&��`����m�Y�:���n"$��zA��&L�r��d?���*�q
CnΈ�b,i��P�w����A�{`xh�).��0Z�vL{���!hXY�z� I�H���uQ;!�t~����F��ul	X�ڶ�<yݞ8=�Cy|����Q�Eu��ќ����yK3���"���8&����;"�>�@0Ӛ����e�����š�g���)�WZ����6��~��^�cؖP���"�!�L 6R��C%�}@���h>v��SD�d�|����d��|V�g���s`9$�<]�O�ӳ�*�Jx�t^�˼r�l�Kƞ�T��i�X�dx��� �ًo�7��|$ajr�;�g0A:;��Y�ani�}ґ7+�;h�/b����a4���ԏ��5K�j�UhyN�D�mQ��^��i�a�(�g��v67�;�����߁?nA�E@�X
�E
޷�����z����a'��G쬔�j���]�u1��� U!�<�D�za����n����ʴ���R$cJ�_v�NC�8��[",{U.�C������&y͏`�=���=��v��!=N�
��N2Xl�C.��OV���pmy����1�6x4k
���͓*�p���d~b�'OgT�ߺ�"��_g6��{�ݐ�?�q�
DL
�~��-�bg,*�F��`n�2��i���R��w��I��AǪ)�������W��G	<�%ӷ��u%K�m�a�9;/�W�o��5��p��v�p�{1`cϑCM�����j��U�����G7��L�����4�D�`]��g��=O�z�gpL/���Z�E�l����
�2���.��+�t'���U'��m4���O樤�$�����i���w��/�����6��.�t�ȣ��`�ڻ+%bK�3�@Y���C>�2-�� �o��q�,�O%�9�D��E��F�H�`�+q�����