��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o ���>ҽ"�p�����6�
f�y������9�#�� B���~�'���Nu���X�<�F��j{�iT�Pv8�����/����A�(�Ȳ��	xq,[�=?[�v��
����)�T �:�zl(dJ���[RTX1�;�U6���U�Q��ߞ<Kůӵ��ȁ�~��[�nV�qΧ�҅���l�9B�F�����������{�IB���[��m���OC��ϰ/4826��58����iԱٞ�h
P=����-z;�'E��ݨ<����_����,���w)S8C&W	�H�`�{n��J�q�oQ&��%:�*#��{��:�sVL�<�O8�9.S>ߌ���x=��m݆�>��	�+�
j^<�I� P��B�^8o��=� ��;d]*�2�0-���p~`�����jC�ЇY�lU�ؽ a�� ĤƇ� J	���>>�a�u\����_^
J8�9GE�KB9㛷筟V*S'5WL�����kr���LrnMOD�|�%��>4Q�������ȩȐ{����g=�n="��x��d��.�|�t����<���vIы��./�!�f�
����i9B����
��E���D�35w�9[��Bl�ka���ղe��ޫJ�w��ҝ��6G�+iq�8q@+܍BKLF���J��z�2�q�Ey),y�9k���n[� 8��l_��������=hNJF�������,]�\�p«���a��9� �"X%PC���ۄ����'�o��g�%s2��-{�X�}NZ�}�j��2���?��X~���_f>7y��zv㯑� l�7D�GH�?%�ʁ�/s�v�$j>��1;�o�MFc"�wyr��O"���TM"7�n����o8'`�/���9��o-n?�Wa�2c�n�B�q��E�[�iu5�QRn�����2B
�ih3"�9 �� X��Ӏ����H ���)�	����q�@L�T�)�Ğ�ҜE�Œ�=���k&�Iy�Ǟp��~��u�RvH��A�J��8���,�%l�>�������x��X>1�]�7ˆo��wQZ�8� ���0��_ �!u:B!��x��>��&��&mö�!q �ұ�;& ���&����iYW��ʔ|��5�ǵ=m�HRꗟ�[W�p^�qb���� �Fyλ_���m9'H��R�Æw�Ǒ���00K�yuT5�t�bG�lzn׎�o�Y�Z�WR��$���e�.;�a?2�v�jֹ�>�j�}Sg`�����1���E�\n�ш��F�Ø�;�4�a�;�>�a!�Hn��Xr�/��FT�>[�]a�:�G�c!?y��n�*?ֵ$�*�`��%�x����"f� vo`�)�Hi �0��\J���|���[�r�"�h2�M�h9��\�ґ����o;�ٝ~�����3Ph_��5����{�4 frL[�>�m�r�ӗ��M51;�]��ٝ�_�F���������T�c���G�葸2�䆵�׾z���D�ѥݛ����Y�ޣ����Iw������d7�*��A:Xm�=|%�d)�AY�N����N̉��/@[�+lԶDDQ��]`ы9�4��(�L����i���9���O�#�[O~��ᵾ;3<���N��D2$V�֢�ڄ��!������f��I��3f�I����7���.�vy
�p���+�M�C�)�ݥ��i?3����Cs��:�MVJ����w�����/��@|r��Ox���e$2��HY��.y��W\Φ��)u�ܻ@��r��z�V]�|�s�
>�H�0TTO�=;,��h��6�ŝ�g��8&^�c�pn����bA�[�ڠ��)|��N�b ��?6�Ѻ�� 2�����b,N� [��S-��D}����d��]�޽��b⯑��MFO�r����!6i5���^�Z�'7�qt�V�9��B<8����9�������Y�î@Ww� ��?�8G��	�Y��
�~|T�H��r����	KL��t�GnR�i$a�g��v  ���>eR�4�dGj��d��PC����̻P�3���2���q9�����^2���L�m�G�ו̂�V����%!�0e�o�$'�����B�0N>��	]��j촨�1�m��ʰ�:13�V�#f{x����"]�� �/�����t]�Λ�V�q���:]���dY��r�o�s�b�ͬ"�����A~�D�h���f��*�QW���>w�x��o_!���3�����_��n�b�G+k���d�n# �t����^L������@I݄uLD��	�L�EL�V��JR����	�dT7=�[���`+�Þ�</A,Q;T��S�����ۯ޻-�/�hקR1��_�_�;S枠�A��K* �z�ځ7N�%��iLuϐ�Ls�����W�f�X�V��{�AHI���ݰOt���x� i��b�^�CGhU{���e��8����K��H^�;6��/�5�fz�*H�T��+��JJ�;@f)G=�J�Z��;6��{Y�7�\*pb)���d�v�pg<i~av$eu�z�\osZ��~���i�GM����3��s۲X^L�����iS�M:*s�e3\vY��Bs�x�D#�	���8����-/���CԃO���g������'
������M��6��K'J<b�s'�+d�k�L�����*mē�9���MO1�)T�7�8|��=�U*}�̜	��'�>�
|������|z��_F��b� �v+ Ty?�E�$�ZH��r�.fm�9�����*wA�o��7<�� �`�R�ǰ�����W��'r��k��TNd�>�-T�B����B�L��YLi���[Q�j8J��y�k�����:��ș��;�{`d[!�~�W�/�\P����S����4\2���ြ�g�)��ݡ1�Mr⩯�Wڢ��b�L�*ŭlS,*&�ׁ�ʃ��<�X)z�-u%�4��#��?t���7�OC�O�����	�{&����4*p���=G=�Ę�=��,b�X	�~��{��7�|��b�-����D��d�vl�g�m[��(.��s�Nce�뾧�(Gc!%��^]��kQ�?�:眽�՞���֩Y^�Q �cp�J����:�w�ނ�k��o�{&4�c(�,�J[��gr%q8sB&[WK6]�?�_W���*��ћK�+�����������95yϥ˙52��ڥ�h�|0Q��̬k�������(1$@�a��x���!m�*�^��(3+K��S��dhaƢ������V���7�۩��r�e���ǘ�����+����J�'k�T)�
�u�A��V���] ��o*��g�أ�T�,����ͮ��9Z��j�J��S��E+��v�ܮ ���[?D,A��G_�9��t� 5?BלLaWҮ,۰�}RW���oi&�B���pG�'��9f���:�H�}]FMḾw��t�vR��Q�?\@ ��N9t�#���:����w����17���J�M�|'��`�w��y�Q��֕�o���TDD����N�Cc�#�dW!ʕx�Լy�_���uR��wW�Ķ����5��Xv�\S�2�I�
�!?'��ʘ�\B|���ғ5��m�>��'^42|���htQ��
��q<$:�7�ME2*Cǩ-.`{n�>�&펾��V�$i��y�Z����j��s�gx�<�+q}�j��=x��1���Xg�@�PkⰮ�'SxTG�� �h^��>�L-
�UƱ�ݬK0�h�����H\˧T� B�&���ʞ\��Y��3�9�*��!��0�bO�i�=N���B�������Y�V\�_満�����2	LՈ�E �6�fCa@��1_�h�x|��	�*$� ~c�4��8�lQ��˨E���d�3��]��p�:�%���G�/c'���@�����_�n=���0����ǭ36ljl��� ԍ��[�pW�Nf%�@���F�(k`jU;)�Z��ޒ�DP�O8n8�t�SX%�7�>����񫪲�L��N[��)��3ݑ����ۙct� ���q�G!9� -U�QggxS-f� ��O�)-�!��z���LUCh��������k�/Sq�[  3���w3#�i߷�)�?L"�����F���pԣ[/ߜa7,�!jr�r��Ľk�e�#O߄��|��oZG��_���G�^������w���u�ξ��[FPA�Ö��^��ǅi
H�������Bdv�������t���H��t�|�Y�$J��;c$���l��n��,�E �\.��^��P���@:�5	;�����&����Ր��y.0�d_�3�����nvjk�.��7���&�j�M�_43Ԏ�ӗ~��d�(kʘ�Y�PD�	l�����ٛ�O��D��X.1��nt�[�i>��hꍍQ�����{�#�T��iN�M��}�����#��}(�BjA�Q�r��S���hm��<vcCJM��a�NL�ڠ縤�4��in6�bn��� ��3�^nz](���U���S�y:�'5�z��-4�g2�3��X��
W���ea���Cl<�o$@-2�$����H��ҿ�U�<5�VK��m�޾;(��a�i�t�	�|W���5_P�-	jƏO���^�$�u���e_��\��.�*+�
/;�0�0��s���	~g�ج��t��=n��#��6�$(B�,@�GKN�"�����߉.�_K�Εq�(���0��N���46�d|���K�;]����v!\��'�%��у�hSD�B�jBa��5�yc���RCT�i�VT�������9�i�"��.j.,I�9�z3k#>�c�I�K��B	S��LL(�/V�ji��@��[��˳Si���\Aۚ���U��Q�mr "���{�?(�GTNeS�5
J������͠P��e�w/m"��-3ܙ?Y�����3)�cP��D����NZ���?D�7�}n�Z�����Y��ss�VMC�N�����>�_i���]3ҏ�B����J5u���js<���"u �	ɷ�s������"������=5���SH�g�C?(uCNL�~;4 �ir3�R4�.}�#{�
��+��IÞ�t� xt�_|��p����Ƿ�w�W�aj-�Ib�����4������&_�OF��{ԉ+<^69���&U���H��f�V���b���^��w����}H��s�,�W����-����ԍr?`�1	�����j��m4�٤�X�<n���ogɻ�,��}i^u����n�!c�ѵ�ԇ�W��oM<y�NYy}�] /*?IW.��O�y�z����D����>x!�Y��c��v�.��Z���QuW���[��k�)_�c�P�7Z RǗ�IBj��]�|�3&�zu�/��N s'!9��1�RA' -��5�����ӛ�l��v�.,�YȪS�����<��d����i�SV����PT?�t%�ݎ������Cd�ɷ�����X�t��i�V�&5�o~?�!�D429�B�%������4&��Ԡ�sJq�����KI`��������6ZJQz�$�JWPخG��������x�r��.wr���*��Z
����Y�h����-S[c��k P��mC�F`pv��s��׈�6�� cf���ʪ�s
���2(��CT�DU:��#��"m}��\{����m�,ȇ����jҹY�qA�SF=��A�7 V����ʫ��Ǟ����e򝝤�Q6�L�	�u��5���1���ޒ���Q��Z	�u��p8J��K5�Y������(s#�m�o<F|�B����R�l�d�Z�����$,zi��|�!A����a� �	�֕_�?��5L$~9��i���Dc�繫�Z����t���*R��%;�����=O�X���2��e�̚D�z�����)�/.�ûªP%L)�&�#[Q)Z��o�Ւf%҃)��;@Xh������N��PR���9 �?��={�������?t�վӶSԔ��"��jw޹���$�N�\gL~����b���9ڲz��g��lα�.Ct~E@`p]w�Tw	�HW�NwB����f ��{���W�7�H���|w��R�M�!��	�O�]!X��@�6ذR�>�n�sZ�؀��޵I�Q��	ؒ�yV�t^�f� �}T���H[�H���2nM�T�t��5UJ��֧��-��?��t{vU&JqA�52r��.t��C��C�`���4�{�����l�B�#���IB0qH��j���]G��F�K��p��:wjY���b��f�a�ͫ_�Y���H鸏�4����u�����JH���GvQ�nt$�A@�rP�$�w�d  ��,��;�7pf�|_E�OV۷�F3S��ƍ1����ٷ�'	��ӱ�.�+YM؍~�^O�\�0���̢�a�BͲ\1�����?�5�zުxmK���N�kOW�1�wϊqd���ٸ��Ȣœ"n��l{ :�!�f�Ļywx��'�����w�'��GT�� jC�s���i���=���.=�X=w�-���/[_��r��)U� ))&�v��h<�>͆�.��W�lM>��������"\(�4g!W.����d*%8
�܊�Z�t�9P�	Bwo0�꾷� ��s�N\��f�o�F	,����q#VU�vo�os>����w����"�6�?~��p$o�����}͚�:N�8f�)�U�a���dǒÚ����*,�/!�IFz����NO���<M�>$(H?�	=�*��g��{X��=B}�W:��\27�	Uu}��6��9�%���]���\���ق78N?�X�#�
�٘s�>J�L]�<�,{^�c�c���Nu?聲����=V��o�hT��3��X��>����`e�h[�A-R�u��6��J�"�)�.��z��b���^P**fM���n�r�D�_&���9�jVD��@ָ�2��t������o�b�H�S U��Y&���*d}s��n�����]j7[j y	�/ �s�~�ׅ��	�W����l�d���i-�0 �
$nݳ��%��v!�˒��%�'9��K��g/�ȧy�)y+y��!P�q��e����-�i>��s�� ��h�X��?�K���2�v7����%nX���\w_&y9b�G�sm��lo���Ћ���W����>o�T{�*�|q��|�6�bD<T�?��$��� X�w��-0�+���п鶆wr�"s���o��s��Gů�/��Azh�¦.fyt}�@}��	���T���u0��*��~�q��r�K�XL �<�ӌ�t�nf�Uo&"b�w"���	�4E&%-
J�U`��P��#���[=	ˀ)�}N�q�M�h;:�{����f�t��#���6�A����eC���9�P��|�(B����ir=c4~j¨��[��N����H�RG�z}C0(ͦ�;��4��[舯��|��fh�S	���v.��.��荃jo�{X[&Yu�j�ĜmB5����^���pI�����of=/�跗ͰPO�SJ��en���(�{d#�	:��^zx\�ϓ��j����^�O��\o�ϝY\p�@�MZ%���]�D8�Db �a���q�>X��I��|��!��ܱ����<!���� {S�S>��5������o�P��<��Z�Q�������Z<����S��w���埔���?q<X�,^m?�&H�����Dظ6�t8�����F��q65���u����D,���EԫΩ�-<�L+|ű�ҭi��Gg]&�z�F�+k=�զ}K�m�fX$��cah�eK��nͻ�&&���k�;�.t=�?ơ4�l�-Y*+#����J�fK�!�ѓH�q�;��n�j.��C��«Wkyq[����N�tL�^|U�B^PN)�c����>5M>�1���r�B/����M�z
�O-Jc��X*q���.�=�f�1�1{��>ruA$��x�ѻ�?�	�kI�$����O3 _����`�V��w��z����5Pi��|��
��l5�#]f��J'�Ft^�U�a�o�Ūf��0�Z/)C�oƶ�c�b�1���
-�Lf�1t�;��靉a���D^�.�/��b��[=T	-��)���M)�1_�DB29��DČo���1���	C�ɶ"�����&&��qq>|����ux�f��a��s)�`>�3�ٲ;P���ոF�g.�N�C�
c<ڧ3q�m�[��IK������ �x?�r5�q~��>�6g��D�?�2/S1b�ȱU��i�\'$��l 0�V�����CVUq�� �e�wT�A0o��A��O?i����X�K�l�D��-����~���[-6��=�/J9�Sֿ�#�T:����3+w_h�+�c~�׿'v��N�7������F9��=?O>	�4�� a"ڣѐ�a]yq/�j��y�G,b2Ģ��?K�hG�VNϺP$i��)]C�����:�@�;����O��E�vQf�$��K_��xtFq�Gye�?ܬ��@Gc���t?��-q�������3��S�ll�ъ�Z<�Y)S�nF$��&�K'J��w�I��tF�ݴf}�׏�V�U�hY���֝�X��� >c�{S=�]�t>K�,�����6�� �g�	�&(���N֒P�Q98��E���%Bc�#�ݘ&4�{K{�D�~ŔѲ�iR+��&N�Τg������K�
Ť��*�|!�M��]d�Ok�q��o��dY.�[��zT˖���Lof��N�P��(�N�}Z�O=�xewV�*��k%e����6]�Q��k��!�@T�E�ȥ��Ћ�9���[��;��z|f����� ���m$E����C��6�� n�3����$�{",Q� e�Z�B�J��;� �c�SUj�UUѡ�O���Tҟ��i��ܘpBmg��$L^Qᬇ)_"d~X�"~��#�G� 8�jm�kz�g,�ݨ	ɲ���b�`S<��n�r�vN!59{��й��B��@��&���	�F�� RJ��y�Wʾ:6H��A�v�]��Ey�S�~�щ�G�u0�En�ڰ��1�ߛҢ�.�F�s�wW/�������EϦX�W�I\;tW.��>l�=i�~��
vE!�!�9�_��j�7*%��Q�,6���`L2�����z��&�2c5�$���� �3Z�Q�İ
Vn�U��XT�&<��t��H������v�j �\Jm;ⶲ��,��Ҡv�	/�[)�P��f� �ռb��'S:Oo�-����8JP	���lh��u�jS����ۓ�L+Z+��ԋkؤ&z���>t����s��Pb�C�ɧ�7V@FL���h�
xtW���rU�_	�wyN�W\L�t[+���o �4�(ʎM�!��Ę+a��V*3�8��/���ۜE6�s8�az�י��-\���  �6F��[UNWr�>��#����i�_��G�)���e���"!�r�� 48D��B9`nVמ(��6�8�둟�`���|3�=�H���z�S@`�3��nG2|��Q�-��rs?�ݑ���������>�+�PV��.�d��r.Eh%�\�O�� ��ʝN�[�+F6�Z2���N��������S����O����e�/����շ�/�U���3H
Sw�Y�L��(�BAoo�)�o��B�~kdrk�n0~/��#Z�,ɰdh=�(����2�VB��<F��"}F>Q�R+ciK`��עHQ�M<X��\�g  �@E�"�g�Q��tA2Y�Bq�_��W�qW��og:�ZNt���}��F r�Lw �i���/A@�r���]�!��X_#kx�w��ٸ�sS�G�z�WSO��ټ��>� T@0��Ax�-��'�,�cdxU1�ԩǳ�I*��[LxqI��Hr��D�_���$�j���l�`�x�@�6�0�O_?�?ݪ���m�
�8�Y�C���)�O���	C�DJ%3��L�H�Bq>ߨ��d�q6�Z��N�CmP �K��V����Gq��1�[}�qN*k��x��Gܽ��a����N��߰�6��'�s��d�k�n?T��Ͻ�p�u�c�ӑ�eKW�2�ӣ����\_��D(��pZ�V)�5�Г3�(�i����V ��P��:�+�p�ib���_�� &i�>���\QO�}�X����^��H7����z�6��yv�3�l��U�y�`���u/�ot�iCq_%�Y�t��ُ��zP� km����+���������y��]gb�����S)n8܎\(+�����9�|(Jc�^�����ߨW���X���۠(��V�f�^���P,ţ�)���MT��n��^�MT�GL�`sz�w�i�g�T�S��saf�+�lt<?K+�쌋�H�{we�_E
~��[�vJ�1I�ʢ���[��Yh�S��y��G�p��?�)r�0 ��j`"Z���	<�C���T�~/�=�$�
���y%�}k�W3
W���Fu`���-��}2�T]����ȿ���NZ�\²�P����ӑ����g�";=[��P�鶗H�Wb^�]w�Wf�4"���Z��:f�c0SƐ3��jn��ډ�3Ǘ�WW6��ۡu#=��p5
����D���8��N���ͥ�IƔ�4�j���(���g��{"|r۠��>���A�VD8�]���Ȕ ge�gQ9��5RX�LԤA����_���2���M�N�k�-@Wb4Z���<m�߬��Nj�7����v:)݁Z�m�Մr���̮�v�қޠ�n=���=r��;��ْ���X�U �h��