��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7���_R����7aPN���BƉG(SѴYۏ~�Y3+�<�&�L������ḍ*���u�6ᓜ?j��{|b-ْ�(��
�����m��<�B>_�$Y�73�^w3ՂR{RC�OS%�$I� m�X�n��0ucj��K��r�˫�}STa�����yy_�]F�3�ڹ�m���:��p�,�����KK��zv�x t���Ӽ����Ƞ��b��Հ+U����v!5�#��01I���K����� �	S�ly�T��Nj�������]bD���_�y��$*{�^�<�a�2㳝s�o�Nf����T���q���&l��4��х�4�Mm��H*fO���;�tP���tM�"�R|B��B�?M��$W�7t+ H�𹇗�SQ��;��
�8vK����(�C1O�0A�m���}i���
I�X�Wƚ�֫d-�����c+ �1u�M�-S���)&�d�H�̕����A|�Qy	w�Ɇ��B�ɱ	��`'%�l����7hug@�m�����y�ݪ|WK���˞��gZ��BK�yo4V�
ɡ�l�d���s)�x��i�Y郈[~���5ȇÁ��e��L���?3E�W���Yw�Rjit�ޛ����F���Nf�>�O,j��H�*����=t�F��uK/~%�F�1�h����9E^K�u�D�|�����R_����s1z��]� Q��$��\�����2Ywlܠ��Sf���{0��X���!�ȎU�Q��.x��@>E�ӑV� Te�t��&|oA1i�c�����b���e���A�DyG"9����!|��f 1�k5� *�1H�����=i���Ys�т#��c�X?Ѣ�X.P �l?=��{5Uy�����ww�T�r�D;lw�q���r��a��;�R�(j�ǐ��y��|�40��7@<����.2�L�%B�dL=^�:�e�LUC^5����"�s�W%-�z�a	��;���_�c�R���R�����ʫA�fƿ#J�����H��mB��i|���Ъ����>/�b����PF�ž�ia!zc6;��S0�~�B��ҝYv�	E�qVY�'�����g��
2�������b�zz�|��^|����R�/g^U�����b���B�5�k�%���y��^�w�-�,oچu��]v�,
�������lԣR1�ΧvH�J��g}�(���H�4������#_vd�����V�|,BO�����0�>���p�
Ģ�V��|�U �o�F!\�:#M�}� ���s3��C��|��9B Ɯ>�mkBޟ \�\��E��'�!V�:*�O����9C��h<~���DYMt�Y�@h�ɣ,$�x24�?W�(ĤS)ڕ|?oH&s˼3��4�P����-�|r���ddW;����Q���D�&�<�H��!=����a��O���`:ʓm?t>-π95a5�F.�F9G�V�"k���c��9� ~h�&�_��|Z�0�Y��8��XD~cJ�۶�<��gHC=���d/� ��B}�`���M�̋�Ϧ)Gs|���A@�1K{�q�NM��h���ĕ�,�'��Ʊ� :����j��E�+^	�a�ZQHxxR��EP0��Y�|Ǌ������IS=�0A���7�[2�u
���2���V/���?�fŒ�I�`��^?�mH�������s͇]IJn�T|Lhሿ�_��B!:%�dL���� �������U�����h�Txf�疹���X�lq
�}�����'4�ǳU*����G�NpD��
�{��B ���;��f�}�':Rf(�]-��>K�[�P���ծJ|O[�u��ܷN.��z�SXK$�5A;�ݓg)���c1�#���z���}v���
Z��ig��p ��i0;|{���C7���N�W��[sS�ޅ�M�T H���zN���%��3�ߦl�"�V��P`lU�`���6Fd2�+y�%N
D<�e�<�2� )�Ѓ�ʻܵ�@�{�O㲾�0,��}�b�p�9���J�ЂM�G��c���c8��8�Pu��D�����XW|��E�dL@L�KVmp�ᒶ55�Fb:%�\,�y�[��U����D�ͨD�嘡�=hL�i���Uk��&ٿn]�8����%�?ˌ��5��
���>R��G>���S�?�Ǹ���8�T�;Ub&�E?;g�5���Vf��g����.�L���OB�Ir�7!6�.K�xn��V�v�WU}^�k�� �I�'I.�Т/i�.O�5��u��6L��q�I	�6���b,��3��0+��^�[w�{�]��tZ�t�v����/ْ�n����28Εj�$�����>߿/-n�5���2��^��5~R7	���. "�$��|b6&�.��Op�����-��v]8���7&�D���I�̄C�l��S�ϋS�x#���h�E4�<悶�,Q��2cd`aU4>�1�t�b�=�J���۸$��R���:;l4tu9`�W��]|�L�a 6�7,��&B.�]ʍ�P%fۢ	���4��c�Ĝ�5�.�4P�����Ύ�We��)D���n�	F��n��Qa�s0}?wvʦh����6�/2ʹ���� �� BN6eɰ�ӎ������a�(ڮ�0N|_p䱜�J��.����C0�h�/N!�3����k� ��1�㭄7-�͓7@W�r���[Qig���\6ʐszp�@�ܲ�s}�0��ʬ��rA��_,�����GcQS'HBĎ�!>��=����#S#$	@�2�'b%#)A7S�S>N8�v��'ͭ4��W�/)U��V���]F_���+:֌�_��G
�'pS������!�:ɘKr�PcU�yw����J�u��¾�9Rz�u���� ���a���+~|�e}�0����`�7�P�l�Wqh뢍���.i�
�ް����N��Y��"59�`��Ŝݑ��F����$�b��K����{Q�f�T�6�m�����f�2o�(��HP����4��E��Sכ)�