��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o娃�dd�;�$.�K����I�§(^ë閤"_%U��:�Ի�?I9R�o<��8dc�C�(��.��`[t�Ƅc�{x�ٸ0î%)��
�1hx�𰳶p��,��n��ȸ~�5 �в5�~Ҕ�F�L����]t���[�Ο����&�=�p������Wu�y73��o��f:��+D���wҼ�J)��$+�DZԤ�+i5=Y��˜L'Ww�7v�Mk�Q�m}�RmJ��]X>k5#�1Ue)���z�Z�0
$��^��4{O���:rv�GMi!�FL����E:��|ك���J ���+~Qq�A�&R�����ц��)��,Ҡ-t�QZi(��U����6���jְ����e��L���f�x�X���v9�o�*�B��]�j
5��y��7{=�N���_��Q��GD�ڒ#��x���a�t_\�P('�Wйx�ۿP����MWDt�f�(2����Hi4��M���,t���t�W�ܻv�Z\fG�!��?jd���!R�v�S�0=��a2���!��D�����1�oBѿ<�#Ĳ����XI��sC����L����������y;����">�8������%̇YA���x�!:+k&���(	�6�]=|��rN����Z-=�6Z�4�+/�����z�5QV:���d���,�����"��F�0	c��H���1*���M��c�F�\��;}�j����$�Hr_����9௯�e<�߉?���O�q����5�`߇��c���Fp8~f:%V�kKޗ���>�� ��E�4Q���9Ew�j<�V� ��<�<��Tix�99�M�ک> 8y,n,�@r{��9ƇM��ɬ����Z0r��6��$�c�3O*�>���&ʩ�S���-���ri[��������T�����Ќd!��b<�&Q�0�u�v|`����Y�;��U��2�Ph(��f�OW��m��ɍ�^<�}�
C���l�aٝv�i�A�7LM[C��"bs�D�T�X6祵ߒf�^�� 7��i�q��?�p~$���w�p|�+u%;U�ۮH\��m�K�苢.9�c�c+H�B#�)8��f�)䚵V���n��xvΔm��y_1IM�k����̭�p��e���y5E3	��Dh�5<��c$�c������
��FV>nW}#��Tc@2�A~+��.��7��i��LK�t���FA���i5����P�HQ���ǑsBwb��K��~������n�N	=�HBO��P���!n)F��VM���ʔQ=_���AM:}/'aT�WU�w��]�pB�0ղ��թM��V��Чq����7%V�ϵ����lF5_iC|�aw��3��P�w�N��mW3���;
��K�a ^�-d����e���{�^�����1���b4�t�	{�ke"Y�(���������Z��q>ۋ�C�����BZ�H���4%�X@����ݤ�t*rFD�k��+h���psT�jV7J3��|�8Ù��2���
j'X���v�LNv�)�� *σe|�R������(�{������t-�sL�ǎCv����`���-���I����hk�L�,&�y5�p��q���?����m���4��k;����U������n�pG�����@�A���m�y��I��!��ɫ̼L���7�eu4*̷�ۼ�̠�GUpB&r���18�ϭ)*�O;�}��M[#-;!�����߅sG��2�̪`���+���]ץ�U�ꞽH)�n�f�|	B��ܖr��V�N�V*�W� ��c�(q�Zei�� ��"ډV#S�(��)� ���*�%gj��V�-�D�)�DHl[|�c�)�i(���A�׉��w�����Z�����L|z�����)3�T�!Ӥ�`ē��i���~�e�A�j�/3>2�#�)8.�,�s�c4������h�n�34�K8A�Ҙ@m����:�4Z�Y�tar],"MRHG�WP0��?�?��H�x�'
���#W�X�$R�H���q�ʝU��w�vȋ>��X�Jq�,��\��^�Q㉨�_�U�6��PM��#�S>�#j��֕�T��wn�X|;X�]��H�tg��u���������&��07��_[���3Rj��������[a�/�\�6MjHKZ��vxٸ�2���=lY����e�8Ƅ�E�z�uޜ���;*F�+l�]�Ȅ%	Kb{��k��S֞7/�V��"1?�0��T�x����pkX���	��'�1�d�g�³��~��O&�L�������G�WjzL�P�d�͛�s=�f)&�/b�~X�|H���[�B��v�8�,��S�e#�{*u����Nr%&&&�|���C����P�׮�6	 �2�<����c�}��R�Mq�$g�c �����j���t�[��Yn��+.��E��i�����2 �gc����!{�@e,�cuo����y�<(��G1�g@s����Ͱ��5����X<��칎�3������:ĶE[�R���X"�kB���Q��O�M7��2����$\f�K���H���Z�m('����/噯*�	&Y���R��4�.}�;Gq추Ai�q��;[Nul���� ���:*Nn�M��_w�������~)Z���`1���J?I�PX �i�y!��E���C�c�}N����,3<�IX��il��}�g�,��W��%���d�<V�y-�m�G�c��U5��D��r2O���_I�_`j
cK��ּ�2�,�Y{�tס
A�O}/��M.|;E�a� �=���u��Q�&ʭ��$QM��}5A3������8=�'���z��%�8͎�Q:2p��[��E��Vz86�i� �9v�S��T�P���5{��J���p.,����9��٠r�w��K��1�V-&]�B	du��SW{m�-+�D������"��HF�w�Ew�y,���ɫ�FdLe�O�$�P�ȗ}����C�Z(Jy9�UY�����uz��h�V(��8	B4z_5���8zً��T�JpÈ��P�;����})����w��o��m��)�io�J�����V2�j�f��>�?��:�#��8��<�Yt�!��Y+����k�� ����a�ʅ��I��U�嫎� �}���Z��P�5�${���u��XC��Є����#^f��-�[!)OO zAt�S�م�{��aќ%���컿(ܬ�;�x.���$��s�j� � ������a���Sݍz)���!�/�����4�L�?��$�k)�2]ip��d���T5��O;�Z��A1R,��d  ���S��G��d�VM�$ν�e��ƀt&�3����!S�%25T���Y�����g^�'�#?�#�Y'�f��9A���o ��7���1�!�SM��T�"��FY'���8Z)�L��/��2�|G����{��а���6,N�2��ߖ�� �I�h��^,����8J�i�^�:h�7&Efe� m�Y[;��� ���/aF[A�ۦ<f�*(((}/����g'�Qv�G��q�V����-(Fs�F�muK��X�v�i0:	�h4�P��:��J_@�ʡٛ���0�x٧mHV�qE�%Lf[�L>ξtѡ&c��;��ڜ�B�# �R�t���؍����GNl��UxbD�dȅzs)���DU/Z�yUrr-���@��i��`Od�����5�u�bI�LK��y���3YF]��#'hY����y�!jn���pM��}D
��PFJ�P����� I�z�2@OH�߉H��1�Y��Q֖f�͗S���-W���}����"��#��֩32�����vJ��l|47��xh��،LO7w�����i)]����x5t��4�!UD��6��PY��>��B����5��7Yp�v��*�z��=y�΅�\�{m��ET�u#M6����0�n����O����T��n˜�릌n�;�M�݈��۩����x^ʠ3=7�y����pE��J��1d.���1:"V�DL �+b�0t�D��;PE�r��r��9��}�8:{2P�����~�hw���Y���-�@�j��)$�ﶢ����8m���D'	'�g!+wAF��D�@dSy)���n���%3	MB��[����(q� @tQ�m�{=�m��&�Br�����QX���y�{�~������@G�.�v�v�m5	�uM����<<L��&$�3�R!���^����bjS\�a��t����7�Y���l}bg��������k}��P�|Ti�,��D�]�/Ou������Y�I��1%�1���� 萲� C����Q_ ,F�e�H`X�1�=�9�卑L>J�v�ƥ���W�;?&�,�y2�6M*n�?�q��z([F ��'��%z)�N@4b����rI��$BD�a6�����N���	���:��]B\���ŗݍ_�F�n�%������� B��/����渿'y��R43m�Zd�p_0����t�<�@������g��Z꟝=�I"NW�����7�7�>�)�~��]֜�s�+�)����P����LLmK%�-^ū��z�N��\��E��/�(��F�T;��D��8�\KD�D�5͑~���n�D@3 ����$�+���E�5�<(S� n[a� ����/P���L)ȖljI�;u��<	���_�P(��!���� 6�E+x9ُ̅52~��ٓku�k2���W�jb{����i��d�j~�#��wAS�d�h$͗D��@@�]�F����w�wk)��Q��ϔ��#NE����I�Rh���.���#\�[���v���8,ɖ�M���c,��]����R�e�A�a#���ę�tl��l�FО 9�H�΅�g��xكҷI�ĭ�����uKY���Q#�����ۺ���o�����CE��l3��y2��`̔�c��%خKb2a�dE�jfT��Q��N���#j=]-��AfYP��|�����7�.C�/�R2�)j"޷�\)�ꇠg͹���D[��bL�['�1fdt���z�9��Ep鏣`�O%@ %z�9`>���߶o��l^BBjj�����S?5hcj4@��{������v��9(�ĺ�6��O�}>�GN�4'��D=�Wn��
���
�t{A�Ms�y~+���ACTC�{N3�&�&=�WDEpV.N�����0��gv3_��؁'���4����:�����K[]��ab�8J"�ZrE��ۜ}ˡw��#����-^��g�f�s��[汩P�#�+��u�l��C�(μ~�VU
M�@0ډ`��j'��ϿP�O��D�����o�,Rn ye�s��2���CP~�����b��)��N>�j�YҌ�g�VI+�5�Ә�Z5_1��f-��#\546���},�
u�[	�X�o\-������h���ǆ�'	F�%��]U�45*�&���h҄��? �W�^���9q�r�
2���S������G���Ї��ޮ﫻�/����	�=Q��K��0��?�j�J���U��ch	��Ǜ;����Lf]U��Qռ��UDhQ�����V����<���wۆ�yU@t7���Z�v@�`��
��E�9@0(����Ë���#��ٖLƚ�ު�K�F6 6��}sF��Y��SY�d݈�0_.��ߔc���?i��_��v��Q/�޻�����ǔJ.�����p�Z�(2�q͘%�J�o*헰��n�O<[9ml}���{gXЫ�L��ʼ�`��I�˙�e|��\�F�̭.%WD�뉵���l,��Q��bܥV��P�}�!Q�͘SOPI/*���<��W�!���XuNi��@o��������Z�<@���	���E�<�����j=��d��-�=�{(�r����&�%b�(P��@r���􈛝4+��p�����-�a��n��:|�� �@��#���h�̛���^�Xs���:񀮫��Q��N�҇�I��P�I03妘�5p�t�����l@H�����9�-�"37�Fʉ��ˬݣ�[X�f)��=s0�$NB6~[x��b�_�b\�6j ۿ�H?����ltR�����<ء�5� ߅���Ʌ�S6P��74��W��V:��� �C'@&��i��w��J�ӟ��5��V(�����k6��,�&#`G��F}�oV�f�r�X4�2tmWg�l�N�EݵJ��﹫���{@`.fYP�Y�i
������Y��}��{G/�	�ɴg�;�O^c�3*��*@�4�̹Ǖ:�`�:O%�f���m���q:n��i"��f7��t4i��j`��*��M�}f�0���)	=�e�LL��#Zг��Ӝ�ot�e]��8�:0B|�C���6�|uI��0'n(��#[Ֆ	�5��]�7Ʒ_`G`�`�Mv�v��)OF�P ZO5]]Xw���1�O? ��_1�ou�tG�A�����L~�C�pp~[K'���"����/1;H�楊O&�m�H54ۭ�M�����d#��^V�q���N�Y�:^�(�O�eG�VN�
���N�&9�A��^o��x�	 �=��*���譪+�u؜��:�7G����l5�<ݿ�|S�X2��%F�_�ar4rG��lQ)��|������N�7#�i�k��
�[��w��Ac�]o��F�bا/�7��BR�����L9��4[�ޓUf��%���`T^9���x5�t(�\�P�1w;Ҿ�����) ����*��4غ���I�����ppq z�\Y�7�����H_�Y��5�(r�b�eF[L��Rb-%M�^7�DA��\CC�t�'�|'FFkn�T��L%A��O0 t�5��mDn��{K��d�ʐ� �����ԃȒ��<g����>� ���=���
:k$LD����R�`����j�
%�1�{�Rc�+Μ�c��.�i�ヤ����_p^����D�I�oҬUB�~!���3>�ˢ�"n�l�9Y�ߵ�l��:E^u�>�<��#Jn?��!1h�z�a���CuҢ9����6\�����e�!5'����3����v���m঺)�A$V���-F�d��06��*d�A"��Sx�x���.����LjD�ѕގ���KS����	�υ|<.�C��'�2�P8�Y
+�)�qDQ �4e@)�څ.1���z�K��pC�</$�
t�C�~�����'�bc���g]{X���Q�sY�7�EP_M&R��=����L�1��M�Ꚏ�ba�J+��=�N������[�Ɓs2����gB:z8���ˬ}3XeE�,m�����;�@,
p�
v��Q��c}}����;r+�ۤު��Eg�0{m�q[��B ��M�H8*NLn�$�:4a�����X4T�w]������8�	��Q� 9��r���Z9$3�T��rxL�Q�H�� A��o~Fq��j	��L��p�|�'���[�e�|�	��F�U4Nz�@b�6���# ��7nk�V�h���z�D�z�
���o[ X�������f�&+�lm���C'�*D�;P�`��`N*/�`��|T3����=8�?N�XUس��5�מ�r��>��%���[�r�
ռ�Ƈ�����7�$�oY�`��ߝ2�+ҟ�y�V��������TE~~����ː�j+ӄ	?�#'H�D��
��X�J��iT�[�m!�x2�g���i������(�ݗ�f
E����-u7�H&�`7$�B�O=��	 C���� ~%�v���(b�B��}��JP���L����"�N���8��\���L������ܐ��Ni ����	ث���cÈ�om5jd�m�9�g%Zz�MT��־����ـ�.���19�T����v�{NQm��$~�|�Wq���z�R���MY�|L3/�R�Y�z�$�n��H�]�K�g����(8�UN\9e�ul��x��`��v �.NNu�$�F��'��~���i/�Z>��S�%����^�����=0.��\�l���B5����"��-�2O�S�E��A����)���5���DN�>U'..��g_�6�������B�$Ff��Ss���*y'���&�z�Ne`��w"'�Y���k!P�����9�n~���ܵ��V0�[z6���,�r����WaL�QN\kPt�Ncc3�
4�F�̆;����2�N	�p.�6"���IB_�簣�Sڑ(rx�-=�%&e>�M��Z���k�Y�&��M�