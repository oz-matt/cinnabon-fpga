-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
A4Y/jCcpQ0uSZPIcFPsPHR9TE7qvl2IFSgHz331tkukzl/gAcEQMZh41JCspiISlbceBWYEExZFo
5+Ahbdl36vFJj+YEPy/1ygaUbG56q6xhsxfikH2BhXKN+7aT62aZxPz3pkwDTJGLIDemCZgv7r0G
IMSer7QsS7vTHdptcQ3mSmXk5mCqFFq8EwAWXBAg39OFGxNqmpS3/+ANe5sgzgawlLrlOnGkkPoO
HapC4/ifeXj4SfZYhAVIn/36l8kqhwJwPXRAwI1bN1fbIWwiYdCVTcBod6IFqEGaBSibnHpXX2OY
e6oTxnxSFF82kG69wJ+IqVs8xWmHFfWDopn7cg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9408)
`protect data_block
iozeI00/IXHKWFc+btXRdOBpPEugzRhIrsgRKHikZQBXncZiW7UMxIEdbjCAxsmakBgrKtlsGxjh
hTA3vnm0hlvLbA6jQzDZxqBuc1woSMiJOlHGFnnw8TDLVuc4LnHP/4nA7AjCZu0WaRdA3MSR51Hc
HEOQut2xhzsZcENj2Q4kN3gBfGgyFioOUYIlXgWaiUIesdlvjE9YKSgDXMXxtu70LYt+nDo5Wp0d
YN+gCL4JO1dwaX9VDWiyimtxCSgDud+2QbYJGk9IYOjW2kqkP/AIk24Z2NIi7EimqlT3PKbv1upC
DtAV7cHrx1Q5sbc4oo2YpPr9RTP2ODMF0qB9rxrhFMji809CbVpDrsLwkSSR/V0RCcsLYM+UOvWa
Twoskig1TO993f4yqVa+fHO7wPcZFM6PsSWPu/k5JeiUFEWXf25POQ7b2R87BQ/YMUJF5jaX8Rl6
ljMw9L+SJ0fagt+CHTHt9zP1Lux47k3CV23tdBWReXa8savhiVYUl6l/bzJgR809/8saIn3F0MPc
2pU36dPXD6U4JawxRNScwHGxyhGASdmc2y1UxA2+BCdkRo9fPkrqJYvtMlP/72kOBLkG7771+AQW
ITwTfGq0Oj50J9Tv7Q+o9AnHQLg97SezBGJ7ciKMKp7oPpmzBA095EmkdnR9nZyJSgbjFtisrgAg
wLjNdWZIAZZoyo55uU8l1Qcs6O1eZPLdN0iigE0R1smjKD7GEFXtatC2YvjC3Jn1GGDd/vQ3FzUq
3/DPXhqw1xvmhXPPnOg3p/WINDkk+gyJi7wKDLCr0jjAIGYozrBTlRYEnDSG7BOb2JLD7jc6sQ9b
vNl9pBDwTtk0ObWKtUNBp5KG42nOZDIlFV8ccs6/V5ZVdLxU20Lr/SfBbdrQNB+OGC2LtAUULspt
2fxv6QR907P7okos4xOhhjUXMnCxYE04ZzTUKSuVep/JvvzfDjpat4oh0kY6kVPpZMU4s+dTGVfx
FkLr2+2aQ2RU7/TX3P0APqiL/bp9TERe2TAfqJUeky3lRHHs3+9WRVKS991bSEsY0Yd/+/Ih+JD2
K9ovkBwcTSVx2AdmsKbY7Psj8JmYpHiSMylMclzDlNUQICK/ZWD4kkqjmdoDULxE79N//o7EJCXz
uoOlJTZrKxi1cUT+rF/h/RtfLzP8bKlcdOpdxJ0cYIf1/CeEcCAUtKdOAGaGYc3F2rbmjwqxLLLB
R42XJrveuGgmFUNRKc6p4maf2eIoGFVoGxab58Db1Y5tBTfunaKbMlZQmAWFbALuZGl5nVT60E3Z
i/4jRin03z+JQcCfFwXqVI7O8JeuKxu3qMM9hiDS/DxW9NCdmpgMfP/ysJbYUMrxaOO37pTnZu0i
4Mc/EvRf7uobY1DmaSoimqx+8BaFGaNTgx4VYBa9kARpWOXPaoe8wsznLVeAhNwGxknwMmNbJQQG
aclnzAhC8L1tuCG5T0zEXPnBr+3Qr8InqneSc1x7E2XvQgtpqoqbgbVMUySZOBAy24ceE+OUuChE
rGehAQ6V1GyJuy9fp85NrRq9WR+BASc/bRuWI9WxzxOjJbtyLPY+ROMqbWDSPDAmTf6LxdrSyJat
4S81qoZ4Oj8SL0fnjHAaSCJPkUy0D7603cKT+DFUD46Wotonr/xb0eofj613hphXuET82VM3IrjZ
hA6dt7fhoGb9mva2dftOACci5dhcwKRcGXFp0MKQFfeSxB7G9MtMEmGHF0hiqaQaUO8s8YhTBUdo
7yk+kZq2mZKrG98bMJtPSR/dVb9gNJu0I1fkIBADBl1e0wHoWByQZ/IZnOcWnXUtKXjcgTmhVOTh
6fr1qtVmWRJX50zBwunRyWDQ01rNQkUb8lh4vkKRvAtL1m5fAoTaMJ9Rd2ZZ4Sob3i1TR9qO/jDY
xQYPYkz2CkHCcziUOkuMt6EJ9QD1MOUcBwGXEwbMlp+JthDtF1r/npmPvcnEgtPD9CJHI6Ebkb1J
xGn7KYH4v5O1rvmiUhTeitMryQjLXGm+idQQ7GoOVzHxeFdPYlguiWqKI4AK1ayknwr5CN2z8YHL
jtZnfFxW4byKTH1SD70drWSL0xx612gHTYIfrU8VW7yBlovqWaSYUL9PhLtSnjbVZ5ma8MtmF3W4
n88DNTFfQz9PnsHEdrPamcUXtzuuFQOLRWPBd+fJFdWbAJp5dzhJIYrqFs0iFG9ZgXZXgXqd9v+G
H5LqaluIranyQk97ciXeRYCNBFFbWiw5dX1we605YB0r/bQ0U9ztYJqYfk6K2NGhyMtjmmwFe1ZF
RlBWkiNVWTzpoapIKjkNz6IskaZ/aEslS0hzhUOuOwmDlqeB1dEHFoOAHwqEUty3qAvRLKw7L5I+
uFENrAEbf6OcJVV0PCYu98pKTwUq6LtV3PMv/92s66sdXb15GkaeyxwUZ6oG7ZJNdhG0Ix8ja5rS
cecYVVny3hH2VPXmjCaERv6gEu56K6i4LLEbbmFJOdQpO0lgeIHo8Ibj1o20yrMmPvTru4pkvwJI
BPaAAYepPvSV1weGbn/bpMvXtHDudXF69aPQfPy9AnkwKk9kcrIwwVzm3Sm5D0rnwL8rqxLTkXP4
ftevW1kpIUnJ3RcSl9DQEEJqmtwCNoQi5/nxoGhs8sbD7OS0hiMnnM7voWgn9UbfPUjnWsSZ4hGM
4kIQCuoAABg+WBBs8YDRJD9rhWrPu/XAwcvTZSb/NfCipSYeDJXJMewMjcgBVL87Hq+syAEeGVgX
0mAtjkpwjfht2pdCz4i1H8wCc/pa0z7+039eqV12IaLHGQi+vPvO0G+JlZwdWn1sRU/1tDlGsqL2
65xqGXQBuVSAbUv6Q0VliX3S+nEKJ9sxve6l20q7iTlwjPTGLQeAO/E5l1KwJNUV/HVO7hbnmyGf
0r4iXXyW13Dye0RSrvETWoTjBklhrGc8ITuCHff1S2X0ocHKFEgTxNYv7ZDzFNgka7gYgEl46ygE
3hUbLYguHZ9Smv0GQgywjK2jPcJ8ESapA9Xm4HP2VC5u2Us7JF9V+QzfFfs2XaL5/0LHHK77OpQx
Ij4gDoa2uufqcFhaThEM86PaU5dug45n7Mx7rTuoFwBb1vYowGveNZOncghqPJ0PGLcFot4EJaTt
9ThXuJWZ45lIwldi33Y8qSRsvk9GbMb6T0qgZbwpGxer4Sd/RtMCKEaWyxME+zPkPTRow1tcecdN
xCoiNaQMcuJEVFO1VbiiAXXG/vcJeby4Kffy8mbQN5XeXUaDeM8t06pSq7WCg0bKY60dTdeNUpnp
fMuiUNmiY4xrhZ5Urijcn5BsJzPo95+J0ZF6GlZp2TPXBICzn/WGdwv1YH17rRpLsVFbiuIKzTsA
2qhsF7ZocI0n+PyTVr1R/wzQ0i8Hax1ZvA/sKKwH++Cs85XVabhnB4Fa42HdI6vwhofDhiZGwM8V
rb3u4KhvKLwiOKpPcK4PnoEvXaOtwKAoGqu8cOXQxpL4BRsIjba7EuDTpsIJjWecpn4L+vpw8+3F
hynP5uEOnMsu3cAL8L36fRgsFXqtuQYwyzOX9rW64LE85Qx8JmAVOBTIzw1866xjdCuFYV8I0zpy
ygbaO2P1EZFsq7SBQ6olEnp4mbh+5y2LI0/kH0Xgn6yTqXLU/bwKozLVI7jIL8brCXJYi762OM7x
6GIrhU7qHrJnTipSGnTREQJbp5n2ENP5IAmr2W5+O/BZEd8gjF4a7GDP81apUUw2lAV/kZXm2SDk
PmE7JY2EddsXEzp2fxcCPHgEEapQoGiebiZCxQr5obyM840G+xin4rVDJXVTit7GRILTrpQteRdh
0JDAZSerw6C7xh0/ycmo8/yA3p8Gv7pzWuKGnNc9u/G/VqwbmLXXk6dAfA3U8i1f4J/4vNBfEfod
Ts8bowxFi5CsGzXnL/vpEwYtQeUKbVb0UlokvIsHhqtS2l8l4LUdkxWTioZbbRRwzI+Xnbw11RgD
XCV7IYlu9pHBcXqDI1NbU76vHTUsC7ftk/P/PJjChkCwi1ZewUQ0OxHCBX/ya8EJPgFOsFSY1BCy
LdPXHDYdH2g6yaSdRhUdFtOVlxMX4iJrXI+H78uWD+alJjEaMjwjivG/Rj+6aUr1pyC+VpzHC4j0
YA0/F3D3SBpk4fwP+3zLwAsBoqTVzRi50F4L4dI6n5i9HlP9d3dOMoVOYAURXJl9J07865KihW1T
6Gde/vzRw3jx5Tx3DKKqWkO+NPBHLJLA93NUTDJMPd6ke0ig2Od+yQ0DkG7n/fW9tWi6XBHjw+3L
Z/2FPKGgQXNOXd23cjLrLCZ7kQYDM4R8U5Zur8ZK8Ik3SbJUp1ns+NNPgl61klnZONNfnKh6eVya
2ZIS+LsOBA4IFmGteveMVsjLuhs+nbbv1vsfCqGWsGn4uu/K2hjJI58M/hZcFkYxGANejz/8znlv
fmWPDSf/o3K+yFlIuiwY2ozHNUVXL5oSpABwZ0Ed4Q0kpKNTnSEbYCxS/V68q3FMy7nPBIc9jzdp
GQ57ACs22+alH3G2E5pWKsAMnAit8lIUqLOdHx7u5jZ0fxCRG8fzcZjRzecb8GOXQDf6+/mHje6H
EnF01wDnZP1fi0sC7cZJ3chdOL7r8oPt49ZkUKS9pfhtDnnr3YAvDHhSYroQYgCpYKopwpmEpYh8
pw8QBlfMNNtqLHtHdsfJCtutqNrYATFOE4rXKhVCDgGtvsyfezo9OPTQX/Q8T0cfYIFg18CxJ/7t
Xbc0NUNBRb8j9OZMYYM4OkrFAd1ooDTqQyCEZiu6qqJVXuhgBaWJipEBzwUL9388TaK3U7Sn7uLg
MAZzL/nLcXlIUXwPCooiJ9CXX5EAmrXfypFaylu6WyWWN9oXI9JTBbiGEjZJU+2KVSyQZxf84NlP
Rg2bTJb0dLSXxcBYiKxOcrjQ0slBFIg3BmQnGZwji/TRlw7ETZ+dCp25xgcLqxjzhee44PI9YBh9
fqmvKCV8BkLrSxZOuMwDS/VE9jTVM0u+WVKQ4JYwFsBcx3BH7wIKGSIx6oAFU1nwwwyHrYPv8lXT
RRxC7jSUVb+tjQwucrJjinb7tQkYuIQZea2K4I3lMsTmpfMNWaIcaZSkpxSYv4SWoQ0RWx41MB5x
dV+XefWznwNkTicdORMH9wuTOzE8vw72kmCF0Yl9vDq8oZ3cKOM+jl3P6unkGphEm5py9G+KsUd+
NnMibVok0vvBitFrgI+GTGNCZ9nB/GLcwX2dlLXk5vfauVbAc2l36YKnEhCARWMZCrR2VLbMxtGM
cucqmaxXesOzcoyX0gKU6BVrM2/twzZir/pLTNmM5z8vi4LTnD5qQFSD2+2cR2LWYEWPrjmgVsBC
eOnQ/zZZDq+IOt3drC8XLo4mqRcQ+h704Cwgyxsm22bmX6pmoRINOeXAMcyJgZv6m8L9i2K2h/A8
11NsN44zb/KLKTQN5hx4CM8iwXWv3CpqUjXcEIRR33PJkS/nJ4T91QSO3C4N0le8b1dn7AOycHVq
X18iw2nR2FjhxiN65KTfY+FVRh1iKEqIAUBxQ6ZUsmOK2P9dHYE+cZevVJy+ypOnBlFeR82n7jJq
F+KycEPn8QuaozeGwYptyA3t/4YzfHre1GmxaZbIln8HUDBQnCcQmp9qaWgfjOWil9cDunVGrbR8
+rggSathZigq1s0/+iN0d0xpQ3p5/TlDLGJLei4sK86lIximqiiZtVUC3jFuSOhUCsjBvQJgYgY/
UHhvdBxrWmBAaNDtUDXahe433Sk/Vw33/NHOVMr7AJl6b3l2Ut5C9Vvw7t3dmfVaS+QgtPclS3hP
mTBxEX9GhJkpEXyT0KWCzPnn2Q0/sIF0TuwRWH+r4fxQ6KRWaV3gES3G8BH5/+DO9zasNZsLtC3B
EnpzqE3l+pajprObdPQwJt8fTM7UA0bQCaVXwcyPUQvJxnAR/pM9NAwyezKMmzzQ41TZMemHFUhQ
WtVrONGf4xJRJc/oWJNYm+LjKkGONtEByXpXTqoOYMLTsn/EHX7s9n6jA/VaWmWjs0mAUbYltSD5
H33Xu8NJX+6z89EJhugfr9ZTm7/40sjX06Q92ruFpiCqBn08pyrHyrMy2zXx2R5soYczwxHCPjwY
togOlVGMD8r+buBWj4BY8fgcMx8WwA+G5R1E90PlRU5FuBJQ1jINvpzC4Tym0oVdqJPNUJQ4SvPl
2zpJY31z4EwKe7mwa6VK7Di+8IA6qNeTFrq+Aa39iKc9ydrp3zXT3b2gfaaP1gqZZrc2+VdX7wLG
p/VFMwG+zBvFxA8Z+wtwp5+yP0EFAJAC4Hy457QBi33zWGEe+s/Rl5h/YRK7S7PLeQgyzZFSjQ/F
4n1PExA/JbUOwxeJ1c9btbeJy2AXiSeMtTJPILE0r9q24p5x1gyd8RDlpNNpGI5VAvYlJKUTCYfw
QD8QrzsiSNRGmZbezm3hIlXoar0IKMvEnhCZ2eGb/C9sPBWMcgyeuK9Xzoz+sAZ5bUIPWv0jK9hq
mnKciV8PIGINVwJToy2HvTVgEIGjXGaKYCbPjGgeiw7oBuKFFXSQw4tkcjaaU2NNt1ehZ/htkCLw
lTyGGuPTQt8YLzDMJHcz0OzBiynKIcvk1voaqCUFEVa0RdfYzNP92L5jts3NxRvttjgP81grwNw6
BZDYA88CDG4qJrX+q7rAh2IUGOpe2zvOmSroqICBlKbHkHxM0GhVw9sWNeICAxuw9KxzkaAj4TWU
y2I20NdAYIkTt20t3WDS1XvivgyA36OJ6Mij227++hx/9VU41FxPKF9mInKf88ak+wYKS3RaI8hh
up22Qz9Ns+nWYNpCDA0bDB86lX0a5+YdyxqfMhWxoF5pjEZmj15FVbLkqOEMePThoztgwTPtYJNh
CaXX8na3/FhO2ndShGCroucXYWgmLXbgAHGx18y8rLWK6OdxKKzlzlcZGBTa88wToCz9I5vAxXyQ
G9OgoW8kMPNCfofzFZWpdQEiNehJ04r8XkoE1eaoknis476Bv6rWORWr4ZIN7q+c3o2S94xkfAOY
syBVg4vSzNkZUxb6okOUsCcjRIkWgdttctbH6qNNZ39FS++QTQg08DjNmkKjJCzCKQD0Vj8crifn
abGs8SeqKf8eiuKYmwpbsZvOHw3nYXFlG2xI1R5L7TXnujcdqaRasgJT8V5lBADj1kRXDBOjSxdH
T54RDKYjzSDOhnZNfqsnFMdMjuMVfg/OJuDsJgr2x0rJnw5LPRiXmmfIY38RVlURyTNXCo/E2OGf
8XJ6XSYf1AuaxNfQjKm5UCyXNXIzlMBcRqsUAXAfuk6tagq4ukDl9Cssd5OCsqH5RH1HpEg6HDSY
yvHr0THULdiPgMp2GoPgB2G9i+EFcl4tHkcSit1djgyJ7qR/EfnHz6s5CUSl0OPZwTUCSDQvLgE/
0+mVJbyNFboAQkeQidxPCMQvWJrgJYL+0QsnrtUM9VaMwJ2X2fbyJiub8baGCVfDBdjrKxNs2ksV
jqN+2F92OJ6j1pS+LYOiYHk59ZmM6qjAYnFzLrYBLDmXeexYzSQ9T/G7Olc/IjXSFW4FukEP7Tb9
KtK68rEykVzfxk4kZd1NF13mL5TGE5LmUL1ykO4a5+YmwXfMlrvvqVRKj7BgcD/TbspiXiZbyd2N
vSYRwja/jAZww2UtZeYBAW5YRds4QYgNePSno/CijK2UkosSoY0undMSEemwxVEIA7MId46CNDTb
yq0sSud9Vll/p6c68p9vwSM7rwMFbbDHVtjNbjjZAQJBBEztsXi8c1+jovCy72yEeG5DcGjHIGQy
CxV+UT89Zr2AD4to9DRY9GQT97GtDLmYXnVGW3QXrVmFKN1rLuvhYYWHsBxuk32EnhAvCd/5S41i
fZb6cvIspx6zJYK9vkJigFMhhfPUOwRLXCyJHzPv4GbUQnCS/+2AK3PaFCLkaNpwupk270hnWpva
EgLnMYM61oQ3sOYCiw76Dq1U3PNp+raOJRNSqF1stpFDn3pm62FycQWAHxqlXBYg4j1JKgy2DqQ4
Pzkqfw2+w1EJH2bHAJ9K/NX68KWQ9QgNaB74zHm0fZLSBG/Jr7UgVhZZGOylYk6rhK3LHtpLxtWk
v2Rzw9mVDftvnVvU35LbKgzJ3fYhetCMl3HZUr6MCH5P1b+OLMk9xL9qCwMBFd6lRoBJJdc0UG+L
S2uIGdm8NMkBcTzWkKDbDdS98paL3g+JTwfLqw+eedFEK7+sedHlV6bhvwZV0GCExCtqNlFpRsiU
xmmwb3eMOYbzLnOWTUFpvZ1p8yKhy6aVY/47kuRYPIOao0JhaCdCZ3NW4Pi06M84IW2yMZp0HBC5
5r10Z5EDEy7hRA8xLXULnrk9Q+4wTRdWs1fTwTL9V6H85O08XqohhkGqxS88VfnOVNKNKTG3WX2V
CEhjyumip1SIdBUxQ+DDydeK5LyYP32XCLvHb0LnyGh3bVmzJ1zRffRjtPMp8RUsLE9x+z9uCGmj
owxzMYAaLXuO1L3UH6xyOlfh+i1Fg7tmbkX6h6rmmudWyIq3czYhUL36QOmHXM39sfo5u4q2pj4t
wgJokjU2GzmdSTqB/l3Yh+IlC1GkYn6AyN5a/Yar0UCrKG1nvtmE5ckU8eYYKP1d3rtycxrCYJWZ
zasnoX2t0a6KDV1GgYZ7mp6uqcJbUXM0j944efn6opL9435uZcjU7PjGPxcTPQ9tZJeWOr3gqm7/
Lsu/zLwf7vzag7uB2eWhCCtwMgAZWJRegcM3IotmZFYpKVOxYioP9R5fsctKlMcEqhQMqbiC+79e
Vqvif6dT8kDOI67Fbzobhe+nb8s1YRJ+7H8cF9PBVyDprfBCTPl0RcRlMTxcp0YCJ3M/Ows8Gtxo
7sjdLWFr0h69Ht5QiMjdy4ebZrGAX0XWOs35yHidoduVtCec7qTmXQI0/E9HjEAV7ddZLpUCX4rx
hzaKocqeJM5F4/4hmuYsyrCPY8eZpQZNU5xBQUbl1NXCRM4siaexUQlSF35d80EyoNJLi58/0EDN
1/gvcwEVKyzkm5HA21t7pj/32a4KiMxAFeFMc8ZOADmSvUhbnuSInSOjzhynogudcsLV2p9oeEZ0
OOm8OAMaQc2xlM5V6nK3HLCf4qz0inaJ5jUvt8p6nn7XF94KDl2FlXPDLkWbjadkcx4cBtP1I81D
Pu9sTth+Gb6AIKWFFny4zAIzLA5zOj1zGiO0elE10cnYbea/PTxbDqFmI5enwweMLD+JZs1jworU
p/pVBdUNV8pkOW8XaO956z7dTd/etqCxH/RZrvJkn0mZIFHVs74gt2Er6REB94Px0Mu6LrCkuQ0F
9w1k6zXV1iWvXcI53L4XS9cNyg/2ZGHC4GJRU7UTo/DpeCTWdOZEBmIN/XhW4gh9ILVxk+AxeYcy
oHO14fVv+jJijay9bjBx0C7u1KXW/YNyPHHuS1LItx2mw+HfpKFANjP9kbO6dKfme5V3rqxw7dx5
ul3HiX9netS4itKv+Dd0r/PhCjo+pl8b/ByCQ7PxrP31VUbAfQWLrjm6O99i7ifXT7U9tyGS/Zl3
edQuiKuRKPip0OgmVv2Vj0Jt7BkoDyxCNwzWav0AXUxkaHjvORj946IMZzHuPvXWbpMN9xelzW38
A3QQtcpqwyO8Pkn3nE76hFGvqARwCFvn6w50lkbj51XtaE/8SBWGIeCGkUdJArYmE23Oiv6Tedh9
DsicKtOeIE3HJpCubtQ8RY9JdRH52x5X9T6His6ZlNgwnj1ihPNFXqEOnK9rmnmiUuSaDlHUNU5X
uLkvG9cWKlHC9g9P44C16FKmgfqLE1ZVB7Hr9pxJJTYFMpF2vLcFbTPNjC+HnCbUY25uIARjb8Ek
PIc2og3nRC8+DMLtvJ/OlMp26+aXacvx4+opG+BR6afDQJ5xXG2pOrfu7qz0pDO+lT1MPd+iMMSq
Kos8bzX8jCnM/eOpFcvNWxyjzXs1+42ZEIVOxRZGmCjdYpk4QAh6yqpbOZgPwPdpWCWh59OlOBvV
txiQHQbCd4hzfbxhRhVJ7s7xJOLjMMvSO3IdwVhs0k78cOF1g0VgY0wvuOcOYvvdvasgrMRVbFlI
Ng9WJYaLgwmi3LVDLrP88E0bA8XK8PGvG62EQmm+BYzkxLE/mJaf3O570je9lRadFQ9iICPGYr6J
JCA3jPzAoCkJ+UrPjYCd/W8/iRpI58VEPp16A8llqWu61eyI565ZbQJMzHL0fmr+3sxx/YCvv5OJ
dTui+2cOswSCSzx/eKwWgFNMjRB7+v32E1aWKJXkNfKN+3RAVJ/SizndsKLdsF6k4ziBzOassJWN
ahonusE2BTKTi0fByeHxxsEbrpibbvZU7c872zV9h0pvC/56I7pLUENvx4M2ZgryHsrYxOAMpOgt
pSpj7kBnEhm3BNFBUJ+6CmBMYdPtGqkyDY/RphyoMRv0Z1CBvXcZjv+stIa/cVreNF5YN7jUx7hN
j96tmmdKwpXoBbxjkpa9Q1oHTCCT+K/z0EYNdosKCAAD27PEYDfM0FmmikQUSPsgRaG1ExMmOYkC
nWznLX7TwkLMctzXx1t0/a2Rr3vwoem0AH0Y2021cwo9oOw9nbPftGvtjSZsCnCOo25To21BOc4i
Zq6cNZIXGq+nrgtXH+25M1Vig7JrBT4gT1awxjvMhWX9AIap/jodtstBtlFRyYdGwuYuZwGQnlW1
gwMcFx1VhFB6JnSd2e3J9WL5jgmujVF1P9ELPQERT27FXFF5v1FMbkbHkn53OE1CPAnqMZ1czcvj
atIKqQdj9418jx2uCN4qiIrHF8fdBJHDNFaaL8MW0fE2tVW//lI5k6cmxlt21nS9urexYHj9Ap4l
4eW5/FTmi4G+4bdLVTAEV/KJaRP8NQK2Iy0i3HeTuv+64xsOOn5DJ+R5AHX6759ZMDzaIv3h3eop
lXZZOf23UI+Is9Jxpb+5XAefzIXBH7ObRTt0ABJYprQyVHRXeChU7dQoyHaK7wG9gv5ZiP0gCFNp
iYsCPsd28dvNVrLcd6mZaSAJJa2qKBLuyhT2kB1mL/7ZHtdR80KT4aaE7OEX6+olyhz23l2tK1XD
Jc+E4Oo7igeqtKeVcZprLgeWZKgPFg1Nhaq+cX+Ro1zy/ICbXgAXX7jaU8uyum89HqUOcV4quUUV
LZnMm87SyMFJH831T+inoMU6wAMEqdHNyNELEAiTGTpORkLWO7eTT9rh13BKMgq/LQmueqqaCPLk
CAwm2hLxCEibmOYFhefN1Y76jqZZSd0G1LlH1mjTB7xeFb0lls4DkcJHTu9HjPr2HbMs59SP4cs6
E7WGw3ekEPNBNCzBfPMbB+eLn3Yci4iQkS1c2YLOOQXNBAp2ITyVs3/q9rGijuqltSq+bIpBYSbq
1gZppc2dNfGdBsShkwHZLRF83d7TvsuCkCoDlXsRzXkJ6jAEt8g4yk78KFLI7abbG2jIGQvzQC1M
vNZ3wjChL6trWegZANM7f0UlH8OEhUPH55VjaxkmyAsrDRZDFnv0hFgUtod3tjh1avQMCufV4FBi
SOBXZXEsZ+OzhUZEFZvjZInDdWSruXFEJyCaF6D1hpaYJtx/oKBP57Wi1by7YoZgjOGuLUcwq7j6
gl6AuFADbwtC7OBItJGJ7c3SdEE8XDNdlwnr5sMz+yVvLXPzay7tZ2fvtFIzzxcMZ/9VL9NsTg7J
q2NW/7mPsVkIOwRVNwJYFrZpJNZM0dEUCphId9DhXK56fI3a6N8POPCa2gGHATIMD6ULgSYZ9kPI
GfxgOQKXGUtTjZlzWToYdigj3EGS90wVu8goiTtZ8bZ9yJpx2MC2fHKRmQ3Nsgw9IX4gGPrLDk7e
HYMJysAFh90t0oo80h8eAo8pp9/B5gG/NbXePPzaKMFyx799rMmWDNZ/mUSFmQpHmQjUMq0yFpke
jnyfX0srJad44P3vFvO9estQkmkl6rux6dWlGn8FiP8BgIo4QfrQRu+5Uox6jILClrgtoKNIS5mT
TBc9ZLq95vReE92I5l8En68ZuDW5j3MXvVV414hJgCe91CxWEAmukzPhpJlMJNVbRwg6YYBGrPZ0
cPe5W1jzHYrepCHrx+KhcHqvxh3DhE9PZl2CTIj10GLDuf0R1hSQXekKLJf6F+lf1j20XlKwD87M
Mn/h2lHi1bKlB+2R+SWh57hMierHdsxNR+cA7U60D+Ba7XKqs7WtEr4E+QbTUdFAVbhI4MtH55T7
DAYXgXqxvQZq3tbcCUCnS5i5FeqwH/hh28yiU+k2KhFnF0Sh3EL/qziafrvTnrdCzL2n2WJHrZx2
23L1/QHhdv1FIQ6P2znhrsTkIaVqfV3oFVq1QusB6r4ZsWhG+omGDz1sXOFcgxe6ASAmVCipShlx
pTvjcJZd9U2jxaoJdVQyvf609IqGbr2BIZqVy1ltXLNdhM42La9gC2dm1I+y9/SjgPQmNlqLBwbw
crhLajdIAAOTaCsZSeaEB0JI+BIrrs1dBzYNa/sL7q8TxqPzUkT5VNTgLz4UDjAM1GQbwkGhd8jr
xZUMT/9DdE7AdxR4ZqzqAkp8aokd3+WTSnARbMt2LL4RxJxQjP+HpIZ5Q2x7fN3tM6BgEBGTExUF
dHLh
`protect end_protected
