��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&oQ�u�ACY�Q�?/#�3�5 /�R�pW�a2߮C��Q���,��t�����m�^vN ���-�2~�	.E�F3@a�=8a�LTu�"��j�s�B##V�1�el'��k,�a-�٪��T�yY&e���Ě(��d�@�����9��+z�p/p��2F���(��O��A~A��"º���I%L���\1�Y@�D�Y�����e�:��yҢa}/�� �B�[и���a~bFl� �E�1t0��=j�,.Վ���r�f�J���2f�!e~�]�XPS"E��_�D�H��,��7Z&�@�v�tc���̄ڒ��Q>����ӆ3��������'��$���g�ˍ%j�_��/+%�������o����@�������o��_�P�PE��>�oT^��VX��@�36��"���Sٷ�8u���wC���^�\#��I+���]�m�`�㺒���.y:z\��nO�5Wd2d�'���.*0��X4����V_NP��VO��y���OT�Zn��[{�#~8��1G.�2�����AB`�N��\��h*��\�~SRk �:�RN9�0�G�CZ�O9��h��"g-3`��\��PK������[�rdi��9��&���·�:��$QM��]��m/j�`�i!������>Z�Ļ����ga*b5��0iA9=-���"���v:0���y\�SaXf�8{Z'KY��B���	FFv�sw��<�6�������[��ù_�W���S�t �
1׻�:H�݊sBK� ?�.[���$�(|�,��1&���3[u<��|f�mGa5�%NP;���О�\x���7�-�萿N<t]ߝӎ:"� ���h�t�K5λGU��$��6�b�~,������Y3�C�>�{��'�3;%�c
	a|h6����� �#���ƛv6�����A�p�袡�(˟���'*ytM��5C�G�l ���4NF舸\)��is3N�����.��T��r�?�αv��}�$)wo@��//����F��lZ�'��ym�%�r�n��}�НܪUssҬ�u��=õk��K�H�v̧M<�d��VSv��8wN�2� G#��h���֦�2����-���[}-�Vl�x�8� "!�lq�w=��5�R����|Q���Z�	����߱��{���|٢��CM�S^G#B��ʽ�)_w߭�  ���4��ѸO~�H���
�@_��hnI��ʕʼ���C����$l�����MQ�5�5�e��^&D��~���N;r�z�QI��4�c���8��g��(�����%$�F�An���z	��"aT�y q��H>�5j2�� J�Q
{����G�W����E��W�n3�(2\_."#@Ma��f)�� �(F{�E���
��|��5��Ǐ-��0P����K�c�'�C��=��ݏ��lJ�)��x�_y��-0�?�Ԟ����|k�e� Igm�.�]&T��g�˾�}�>�BA���<-��-�����T��2�X�xjZ5�|M�����q��[T:�=9�WC}���H7�s�]�#��MFM�K��T0�r.rƛ��)ף}J)P��m���6������.4Lw��x&X�@*B���_6f}U�;-B��=��1¨v�B�^��	�����}:�!t����$�RB�yc����<{ ��Q��6:�.>� �ӂ5��z�9Y��h��"��ɟL!ڌ��7�xr�;���ʶ�S��\����G�@�jvfګf�5�����U�#?�$]#j���{kq�Oag�$�@���|�CF{��%��Y�ލS#fݟ���� ��fu��9'ł����9Hsw��>'��M�p�����f�p]��"}8؛F�Ph<�6��s�#ݱdG<�s���� h���{�֮2d�/
G�7dJ�S�����ݙ��Mٴ@ �8���;�T�>	�
�u��
I󌉵²��-��%0Mvz{b�����Q����Le�^ު%1�}�,;��.��a-2!6�y����[#�-5XT���+�����'����$�פ������������	��1$����-�k׀�%<�y�Ϗ^M��}aE+�!�*הB���IT��kI�5�?�ܣkγh�M���Z|H��>q�@/A��c�+����P��9��u�}��vJe]��'�տQ�S4���ޢ@J���` �H��=���z0�wуѧi'4t���@5�f�l(�W��voE���������O�_{���B�5߳[�����o��OH6�L�ˬԕm��qN�p�Iz=b��n���c�cZ;#Y�["=*����6%T�g�5�J���ݢ��OV}�	�f��B�~<(�������c����R
�6����X��%�^Qb�D���[z݉A}z)��qD�<����a���m�,�F�#h	��`+��x8��?x��� �iFê"��_;�4��(Y���`V��mk����+��B��z�V{�Z
��HJ���.1#3>����ǻH}�-�!װ�q\U
B~Z��V.v�D�*E�J�J\�u�GChB�JS1���J��3�M�����!��q̧��L��OtG0s
]�Y�j�h�^���/�0�Z�c�h=��T2�X��ޮlW'?�t	���o� �:2a�d]�Z8��1���S6���4#Df5_�r�� p�.��'t�n�I��'�Vό?���A<@��l��r5ԫĴ�
��� �,��&�8}+LuC��.�6���Cu�pf���P�U5��RAT���J�9\�?Y��HS,����a��眱I���u� S'�`�!w�[Ue��0s�oÓ�!mѪ�A�(��ٓb)��d-�Q0ll߃��	��6W������Dw��O���~!�?��������S�i�T�G�����o7SQ~𒚳�:�^�杖CΫ�X����QY%���u�K�"B���������1���&�q�!�i�I�XO5�[�8IBȤ	�F:�d.�_M�����4 �ܥ�����@�F.1-c��H��T��8j�ݸ�;o��%�C�$?�$�r9�!'�o�p�`!u�Fv�j�%'4u����K�~��L���}��
��b���a�fXӸnl2t!�4��;;v�Ϝ� ��;@��y����a�&h����31+ �?�����w�R�I:�):I��i?��s�;������	r\uP�Ɓ}�]~B 9It�r_��W������QFI#v��Ͽ���������#���)yyB�)艬�cx��0鹍^f�J�"����(���h����嚱�;,��;�6���PP�Xm�P6�<�
�*T�J�|Ġݮ^|m4�pTLu���Fc����g�y��s�G.���4�lD!EXX�,گ0G`!)��*83�O)<��C��y�Ze͂_�W� *���"2/��֯>k_e��<
ŗ:I�ӎ�f��64�?^���$Z�FTc1��&)���\�bq�=���ȭC! �7�:�2�ա1 Вze|�}�曰�5�>�t�)Js�-x\C�Z	
HwC�zmT@����8���P|zK?ᅜ-K��������Z��S���B�HH�Jte�Ii$�Q��8H�p�?�X�-̐2���T4��� ���]�1=~Ċ$�6�ak]�����{0��>��,^��;�AQ�tk~����<�x�n�
��}�\�޿n���Y�s��o�	��#����I�h9b ;��)y}�P�t�GQ�=�V�L� ���4F��g�A��戫�[Q��M��d!�'	�����MH��T�[�IjěRhst�b����Eq�=A�����
��+�Z�d�%{'?���~ ��3:yT�v���6�PӸ,�:�]H��@�j����|��\��Y���1}�Eba�f#<�87�:���#�v-��B!]B�@d�4 :A������ù1S�ӭ/d{��*l�88ok���~02VʿBH��_4U��!�}��w��y����n%����Bx�r��
]����~�j�ű4��ydr��~J����#����]���O:'_�_O��r\Z�1�iW��<{,��0;��rX���Ja=�[�T��s��l;ܲe4J*��2��de��_IU:`�I*�"Z;B�$��T�b䪻1� `����E{�y��=���V,_�)�e�*_{�gnK �U�'��N��[~1t���u�Y�;����u4�5�5ٝ������sTK������k�#��37��!c�X/�c����m�X��o�F�׶�C�^� �ȇ^ 6�y����+5�z3(�|2���y!���8?�0��҅�`�D.�� o�V+_�{yQ���hQ�m�I��@H�ޚ�$K*V�B�X%�l1������5��I��\�K�o#H�qo�5�
_���љ��ҥ�5`�;���Y����P0�\����U�k׈��H���P�'�d�0V���枫i�Dw2sIdt��~S�VƝ9.n6����֯;CQP+�/#.�-��岞b���]B��O����KbyܒvdDLx!�-��(�^�Z�*(�Q��Jp��Q�_�r��}ehT���\{��{Kbu��$�Y�:��[�I�i󏷖�vo�6��Xˆ��jb�՟@@�f�$T?x�kS�m_�Z;�0%=t2�X�����
З�^���~�^��ݯ
��7�*��1�o��>~lλI'q��Da���[�]T=\5r�{�=�]+���N�sH"/ܸ�=Ze:��u��@)��N�>����
fG�Q[*���q���]c�ݬ1:�?�4���:zR��G��a]���oZ�����-*��߫o���hn| :�w)�<�[�_�Դ�3��b�4� ����j6�~v�x}q?p�·�DIu�HON�2;�r�02�.�$�O?쥙,�R 3�(�#iƺ�� ���^��	.��_��y)���R��˂�%�4��V���ڑó$_�%W@��4��U�e\\��npi���.T!vK�H���$��.��_��N������e/�zF�� 4�<I���d�����zHω����K�j��E0����Iw��G@�ψ�_����я]���e��=M���xS��)���_��2�E��?�H��� �����y>B\��C@�Bpn�{f�ۥc�n`h�7�,���=}��`��NmG#��k���}w�Ad�����8X�'iFl[,��X}�~��s�ʬ�%����v�8XY3�),�Bq�Kn���1u���Vک�B������曌��k�1\�q%ՠ�h��֗P� 8�GtJ���[+�?I��Ap��~���.
QĔA4V�D?�i{ڋ�]��MH���Tjߊ��፥~��L�����6M<��i�'��[	�w�cj�w.1���8 �C��&,��Z�+�]9 �(}iq�P*�=�@�'����'�`ӧ��X���J�%s���𶲆�j"_S�vPf��`J9��V����~���o6���4�e7�5�T��e�����p08�������n��t�Q�(NX�������pz�G���ziM���-�c��Gl�t���/\�7���C�5�:� ɠ��)�͡�U@;���r`�xb��D�i�������go�״P�I���i���]��j4g�q��<�H>��.�H�ӌ��Л�y��'�(�v��m���O�[��6�G��,�#3纣!;ٓ�Tb��qrlC 6��[:>B>s�NUx�6�xm��Ҡխy�W���������>+����3��2)da��~��
�6�� R`�ov��m2�U�!�E'��3�Qu��銯���j4by�>��'��"�Ow���U��h�x�(�_!�V9�y���2?o�[ͪaU	{�o7����P�����͎=c�C�p)5e3��E�Bc�eĞ��&�Q�J[}�=[�kD"�
@�����"A*�#��7�'䍤�BYF���<.��m%���S'o�T[������^�N��x�H���x2'>g*"�k\�Covt�-!x�o%1�-[*9�E:�5�"��^�,'�<���22�y[�2 QpC�.e�����Z1�U|cF�y�/i�H��R�m,�e^��$�SN°�h��(d��W���"p��ZA*NyO�}r$Y��w>�N�|+��☶C�SR/+�I�5�=�>n�l܆��2{�
��Wz}�
F�N!�� =��M9�K�ރ#K0{���u.:Vli{�K{G�i"�q=g�m�0�"#�r�]D���A�4�.?�fAǰW��{_]^w�-QD�6mqa>��#Ն�l�(������M�<& ��=��ŗߚm����ϑ����d��������#y����G���Fb�6���F1�/CU�#�iǶ�\��u�ys �g�������ʹ^���-��iA��{�7�|�L9L�
��5c{7����
�� �@bNT��U�[�ң���0��
h�H�3% �e�1��L/1L|#jڃ��\�ة��Q�¿#y�����(4D$hn�`�
0Y����꫼q�\���j{WI8��詂���$���J���[#%sD5sRXh�,����6-����5ϔ���?%z.!q��͘ �4������{���O�9ܗ�>t�!��!�[�U��
W���"�h���IDh��Ks)NZ�Ν�����3fVFX@����6���׸VT����%�0����T`XW�KI�(t<�f���H��s��Q���;���a�>�����_��r��w/t�$�G��b�����Jc�=!0��!5G!n}������x�T��{á�A�ޖ�7�S�w�s��d�������%�V�{3�$ 8�}Γ������8+v�Hc�7Ӝ&�uyْŦt��?E���Fァ?��`APq�^|���@x8�>���4��rO'3Y�Uʟl]����P�[�q]��cP$�����	4T*����b�c:~j_�Ήڋm�[��l֒��C�UFp�`P m�HiJ0�5i��V�{`�ass��;s_Y����7���cL.�ϘY<��ֿ�3+�.�Dٞ�I��g��6�����&J�$��f#ca�V��5c�̶�z	��|��k�ʨ�6.`a�o�ڐ𤍽�t�F�bC�����sgУ�K�b�%�����Џ9W�Օ��5f��LEqe�*5�|��D�$Z�jC��}Sŧ.�BVh&�xLz���!U]�����������y�F����By���-����'�ǃ��'��2�SE<���8EL�.	k�;��p�D��R���,�vќGŁ�%\BUMy-��ԕ3�{��K��U)�$�=2�/��|ޒ�Ƭ�{��g�[� {$x���iQ�^oN�C��9X0ŭ���еh��L��^�2��q&�n(QI�XD�Q��υ����6d1�?2f�q��GP��� N �_7�~�\y�g~_!)����n�R�z���E߳�jD��3�{ ���M�S"i�b`g�f��8m䯂�v����Ż9b �&�O-{���`�C av��/�]��e���%tT�Z-��o�6�aDIp��-O��G�.V�C���w���S�#�����h�@�ҡ�@���V����0-���b�x�J�M4�y��|;��h�{K��U��@���eH�/���� �P�3yā@�5ɿ�f��4k硬���P�́������ڱ4��ﱿ*��+Y�c�9��:2�H�Q����Z,5�yg��+k��\*U��_6m�d�O���m��7�6�� 	�Y<٦�w��=�CI.�ygxL�
�$�ɤ]I�4����-�^|R;5י��E��Uz�����M P�|s��
���XS©�C��a�\S"*Ma��1m-��(�Mo� 2��c��۫�Kglף[)��E���_!�q�N�faP���BS����Q���]X���yr}|�V���g���������ճ�Z�}��cK��X�oGo8�rA�`���"9�@1\	��J~b@�Q�9̀��~�W�y�7K���	ީ�:����������%@�Q�nJ4��pe䮏�5V*JM��:��1��\r!05"����A���"k� ��m�})��Zbt��(}t�&�a��xT��	� 2����y���'ͣ�3�_�Q Y?�ѐ~+%��uÉ�p����ǳFi�I�4��!X���T�\V?�*��W޵
.D�T7M��uj8��p%"ceثH��f���g����56؁I��6�j���fx��T�_Q'_Z�:�ב��k��8�ֿ��z}S�c�RB�mW~��K?�qĊG]��V���k��A�m��	u��X�Z	�*sF�Lǣ_{&�1���! 3n����(�c������(�&mK��`�8��8�$���J�<t3ڱz��?���d.!T��/���q�;��$.Y�A����P�p��Ƹ�$�Փ��K5+}8�B�L�;��^�+s-�.���L�FD˝��Jq'|�\��^��]�Cs����C�᳙�֕`��O�cߛ7x�굎P �ֆ�byN�,sB��ZVf��$:��l�CydI����:��!����
�����Ȁ	��ۻR���O�0]X�܇��w�{jDm��-�?4wA+c�:Z�G,���9<��m���*�tN�Q��O����"�W��a��W��d%�Ћ��|'U�-�n矱
�G�ƣ�I��M����N���?�>/-%qׁ뚏5�iE�f1�U�U���;��������O�����5W�F�}��ɼv�_+�����hV���B/�(�|���x�$ε�F.D���1ryV����f�|���ua�@�w8Nk��&��,}M����V��Rk�S��k��=�Yt��6	�5i{B�)�4G�A��nQ4΍%	e�L"�����h)�2�̠��g�\"��p�z�1�.�F� k¿j�%�	-�N�+Q�����+W�>�XF3�8[N�[��w���s�e����V��1�!S�%Bछ�C�>
붙��w܎�'QΐT�B�g\ud(����\��g������J��)3wCw��
!�n�����U�J	TP����5/=�&�[�W��.�U  J2m��3����D�����_���<N��+��慤aQ;��&r��K��g��o��mu��C0q1T-�\�)����թ�&FH%����b�5�I��Ru�"��>?3�P3�[(�����,����9�!߮Q|�����"
3�-wd9'�t�N1+U��*�Q;����,>�T�O����K��%Z"�~���,���l�� fr��a��<���Et${֤��JƾBYn�E��g��f	 ~����JIk��"a�A��3M� ���`U�����~���O��t����I1l�<9�[ɏ�����]�Mwy'�y�z1�����Pj5"�F}H<\]�(�s�`��m�6����1��µ|�B�3(~���b�n�G�J�K��G�w5��A�!�]'kh+�#�\�d�G��&�[����u������8&7�3=/�����k����E��KձJB�	�\|�dL^������t�x?2��C� q�{���q�̻0c��2�xEç���n�v�P���藃��z�#��,�����x�>��[���j���-�J�NiTGX���:|H�W�`�+�S��y���qP��O�ݘ�z!k��<�i�w�D�K3-I�F,��/�6�9]��sm�[���'��1$��³.�̕aM����C�\s9��R�Йbȶ%ϟ�K�O�̵AL>��9 �ޱ)����]6D@z_���a��3�<��/>�=[Qc9�kГ�&�j��5�%y�ٻvͨ3%�֯!/.~ی�5s	;�������o�yoP� �0����U�^�w�ݔO���hP-�ե���-|��7~eT&�]���pH�}mb<����*$a8����xX�;������υ���V�$4����q~��|Ya=+�J#%�����Fa�p��L8�Smޒw �W`�~ �K�7�{�q��^��oy�0W��$+o����х�VB����xm��Lm�'�z��B�2��J�<~�&���z�Q'���06*G�2��r�漢�?*�r���>��'��l��d�!�GWi%Pŋo��~�kl���/1
�=n�N�N\D���	u���0h,C��$˓�i��G�(V|�-�|Mg*aTz���As��i��0�;RD��+[T�"�ql�d%�8y��H��|�^�y���,��t�,