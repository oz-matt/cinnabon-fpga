��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o��a�cmU-.��-��<jC���88���i������?6���k ��E�l)A"!j��@S� �F���I��t��]�z-*@C��{{�ٽ�LV��/,�}�e�>>����\���4�98�3Δ'�������Lm�y�QrZ}�|���e U�f�W���N����kw_� �c�R��b��g��i@T1�T5�"��+�~�l���~�B��i�Ξ��a�d;���Ql1����:$�����m\�}7��~4W���-ed"|�Mw|�Y�N"4�F��α
�n�)�Sp̏@΄3�$cΌo�\˖n���b���P��nkO*��q��_�M�[�+c1Ÿ>1��/w�0Z;��Q�� /���e)3_�^���?ģJ�%O���YT|o�ȯ��X'Q܎���n�/`e�G��{Ղ�]��ֲ0�G ��etY�3�\�}�P��dO+1�u@�ؐߴA�7��|�Ž�\��Z�v���{������?�}�X����?˦I��WoU'�>�>�;�*'�G�H�reVXJ���6y���ԫ�|D��ԇyY*,j�e���~;�����e"bלo�|�S��4��}iu���[�`[�� �	�G��0���Pٍ��X��=*J��Bh��PO�F�v�W��h<@ڇ�I3�����,��6/Ӧ��z]�M��w���I�z��^%����y�(�q91�w����tN��m1�42��J_����&�H�إ��1��A��Y�-�)����*�).�u(�7�H��W�k�%a�<;%+�5���S��&2�r�f>Lr~i9W]��;B���vׇ���{ϡf&�?ZB�]?��DzMA��6~�*dƚ}A�'�F�D��}G0)����~�W���ug�Ҡ֧�G��Fm8؏/��Ov���T�V����˗�i�墳��y$%��
�$�g� ��\o��v��Kd�a>�!Զ$� ,FDA������<�VȎ`툼T��ߎ���'ȭ.#���b���V���S����u�i��E��>/�>r�{�<��d��D��}Q�b0s��:h�%c����ovd�#�S�B^��Y�P i�	��7�a������A^�bȈj]������R��{�r��>�2�}���Se�_��yW�V����E��� �:���Q}��5�y�#ra��Jz'��.��>��1�e�;�V9�8�6B�Nı�������܈oKx�zܶ{E����Q���f�H@[�������ǩ�c?����ߎ���\`��[�.��;f�	*.$��<#�<�E��	���+7Q�F�#=���[{̙j�$��Cf`��~��}ʽ��pP�c��ʙ_�Cv�l(b���� ���#�z�̨7>�+���b*���3����r��yO������F�M��Y�B��$S*) ,~\�{l�M����_�w@�����Qw�^�?���ן<Ȓi�6��w-��<*�0n���p!l�0�C'��*g�� �ߛ_o�'U���;fe�wFu�k�2P���t,R35{W��R��'����Z�t]�S\H�:iq���̰�8U��<2S¡Sќ|߇�5���L��p����knKM"�������"���ԟZ�d�"���?V����� �=�c����ִR����0 ��aԂ~���Κ��X����Id��sF�+%�̀�[V;Ǥzw�Y�����:�7����|=�=�׽F0�*Ft�Z#�����'wH5��=lե�;&�
D,󏐟�v?�d�)8��U�k�pC,l��[�k���/����NB)�g�&�\g#�����iF3�-Dhs70�U�;���bA�x<�7l{8l�ͣB���1]�����x��h��BJ�E
^o՛vz���ɚU=�$	PَV�����yŖ3��ì�3�^�^<�62~�Lt�r���.�R�y���tM�O���*{�K慆,�|hU��=��ڬ܎w�>�(u�3@HܾȖ���	�'Z.�9����H��F�{��1�����>DO�q����h��w�&��c��Vd<��*�y�j�.�";�a�l�"ٷMA�N1`�ޢ紅���Oڅ�-��ZF#���6bݠY��!I�CB�␻C����)�$Y���G�r�>�ߔ�h%�r
�(���[��f�e��x�B�(��30qI%d������E�0���|as�W��Q'��bS|��k؋�}��7O1:Z��Q~�;PP�65GZftBRBǠ��t�JF#��ܚ@Zs����}��*1	�Aߪ)Ȯ)	��B%�!�d���л��lh_�x���Q.����S �ogC�k��X��V]u��
�ܳ�.��g=�u[�ӌ��jN�
~ʛ�O�!�j}� ���`YCc�,�ܢ�s���H�hF30��������1�9�?1{�
��+��6#'\�Xքq���t�,��2y�P�*�x�3�^��U�C�4J�L> ɣ�
�����\��(κ-����l���:2�SO�2k-�G(�q����5s>���X+�(W6��(N'�n�
���ˮ5d5�!���A�/im���;��m`~����V��D���ͱn��u�5u<�ʹ�p}h`� l�_
�D��5;,S��X7����c�my�i<9w�2�S�x������췬<��բu��'FgRD����� ��0���~�y�ed	��_���8i�#��>�D�AگBv���7�.G_�oͶ!J�Z:Ǻ)w��Q���O?��d�������IC$ܿ *TW���Ƌ3��b��Za������K:Ism6���=&ھ����7����k�~��e���ࡤ���fn��6�"�����:�k)�G`[d�1����\���'�h�:��&����A�e���d/\�Ƥ�4����4�p#��Mɺg����#*� f����(�{ӕ��w׵�iS�I��!Ut� ���ڨ����9%M���f&�Ba��FqhG�d̅�f2]���z�ᆓ,N(���%2��)GQ�x��[p<�Bͫ�қ��*���mj7��/A����<~�s���|�V�q�=|�r�ðI��dw6��)��ۣ��~:���=�>�����̟S\$����׈���w+������=o�P��/��)*J�ȴC��3����Üf���] ���	�Q���J��R[I��c�K|���&���&\�y�B���9A�X���.d�5�l�E�;���w�:s�l�H��thP�N�;�ǧG/�m��W���S3�$��;�WyC�3�q)��!��x��xkZ������>��N}(0n;Hw���g�/P(��9f�E��~�W��(2� �m_����&M#�j>�γ��*?�j�s�S��E��^��`E�h�C��&�£�\�(���s�h�y�6�=�bZ5��^��>�'B�ʀ�+�%P�Kh�ϭ����
���q^�i?K����uyҔ~�;9�Ǥi�ٶ~G�:G�R����D�V�ZBkA��`��?3d��e)Z
�BJs��f��.;KMyb�] �)�	�x0��;�$�ć˵.��^�0���t?�[نe[�	���y�7��|N��WA��mm9��v �T���Bu�ۤ���(���|�y���"eU/����k�B�u.�<���ds��{�;�+�_����a����Ƅ��E�E���ѣ �$�_{s�8 �8�ؿ�iG���L�Ν��nO�5Y�m-�AF�3��8��H��r@�d�8&�-�7��)�<�%�r�	-w���tL9�� ��g\�L0|/ٻK,Q���ۛ��=6T&���}\��L[}��q�\���8�d��:��s#� �*��k �@I�v�_JV?��;W�b� � ��h���\ZB���`�'��?���~�Iy�j>���4k̓���w'���b��\����:_�Nk�`��,�+��'�6����ko����R#?J�/�O�GېL��&���?��)�q�s�F���=BQ�~�J�]�M"�*'ҩ4k��!��@Sg��{Ab��T�~잚&��d���֋C�7����7��h9�2�ܘ=/3G ��Fexq9ܿ��dZ�c���4%5��u+jc��ɜ�'f��#��E�����L�ܐ���I�3I���Fp~T��g+�D�h��̫Zc`���<�����;*-��ñ(��9�> 0��#V���n�zzo�W�2����gL��{ m`k�MIc~�\�ս�ʟg�L���/�����1�퀬�=��.$d���I�
�&hb=|f�`n��j��F�o�9ʐ��]�2`��3���Գ����I���Z�=�q�#��Q�Qvƀ5��V��(�?�s=�m�iT���Q�؃V_Sΐ��5�jFHCF.�s�T]Z4q!���>>�s�XVɢL�@��h�7�9��2"�a�ٕ��[�ߏ�+d�/@v([)��b_�/�)��S])?9ܱ��]X�xM)t@s}�Bpn�
+)%_�P%�놋��>��_�)�pY�vk�%��/Ϗ*��E�����W4�`�¼�Tڟ�z��%v���p�A����!\�P��C�4gY_�g�a�c�Y9Fs:T�EK�Q�3+t�
�EE�d=D��/ �tU�ؗ�{�K��M���ݿ����蠕^�SK��� �Lk����$Tl\�"P�q�����0y*R���-*��}����k���V.���Z�O@��&T���r�7�gv�wOF��r�S��`g0SPL�<k`�����ۙn.��4�2JO��c�'U�T=�'Xz6���*����)t����r*qN/��p@�0z�>��J]j�#�/�T"T�E�h��I�y`[�X�qt-?�F�����]�!?4Y7[�����b Y1]�-'�K>rf$�
%b}�uDʊ�a����
�&�2�������]�X�th����	��Y��4���~>� ��T�`.c1�	���Q����Ak��yf_��Yݭk�2��9r2�}�$˕0n���5��R@�ɖcǏt>y'#�N���i���,�Ɓj�goB l:1��_,�@�IObsv�'O�����$�SMҦ�œggr�eo��rʈ�xj���uQ�I�b$Y���	|�Zo���)!�T-��KZ��Z7}E�����N�!�L�S"W�-�ɞ�2'G e�*o;Ό���7h�n��-����҈QYQ>#�G���l��1�j�~�����o�QVn�]u���1�hgH�R�QL����o�x����΄�9�'�A'��9�	��WMi:���Z��Qz}et�}#^�p�r��s�MԜC#܍�uf��l��
Ƃli��7���Ϸ%��.�}������QE,�
�����
w{��䌕�1�UQ��g1]Cj�!�v�;=��YBN����\}��)SN�X�QmtĎ�{�˕�{��4w�RB���fi�x�����1�Dȅ�p���	�D7#�����7�=�����$4�3�^���5X �Y�?0���0��C]��f��u�*؇<��t�.ǣQd9O�$��A:�6[b��(�غ����AN�c�3�>_��*�bM̻O91�gY�c<���<�m(�����#,�{|�.Wu�$h��J���,1�|��:  ��D�
�����x�7L�Q~�����K�cM��M�̾ZɎF�𫌷	+��f���p1�A^8>s�3yb�6S��{u��ͷ����ry�=���1�',�H"���誊�>]<,�&�[R/M'8���S̴��\�*��һ��������/ȓ*��GK�%uBH�La{=�<���d~Co��ϳ3؛�L��M?Ȁ\2�	���o�_7��+��<h�rH��4�@�s��m0`�=~���K� To~tM���\5�O=���/P���ˈ�Ӻ�blc:�Xް�6����xG�Z]yW�x�o<�{.!���~�~�� �9�>�7�K~�6�+���p�[�h�,�OU�}xM�&�<���6\x��]�|�
��C���Bf_���/���?G�3�%D�K�\l���w
���͚�S{Q��vg���*�d
Q;���6��j�7�~J�P���݅�:��}}��y���X�����2]s�n'��|u�eP����^�t@��H�bF�綸�����쇑ݕ=7u���[�X?��M�^WdMù�����CLEJ�+��lY�g�9<N��#��W��۰���^ZU����\�Dk�	t�i_���Hr!�.��j��U�]0�l�.P��+RbE��ٛ�	�&��Zp�҄1dE�{�|���KUݭ��<�}-5�.M̠;�9�1&z,���1mКdy��Z�'�T	�Y@��!�/煰�#4{��;h���Ϊ���i���SfXh��I(S�}HL������t��7�G������nXĜ!2{�Y����<����A��v]�	0�:��5�3�or$K��^��e�<�]ΐ�1�؏_�v���"��p�}�i�*��l�>����2����ډX��78��H���a���v�V�"t��[�Y��3o��Ҿ�����V�:TI৅WK��V��]-����U�ƚ�	��	�&�J��2,�`�����d<����S�$����Z05}xkc�h��~���;u<Mo�v��4�%KJ˫)i�+����!׼@�h00�r�0&¹8V�G>݆�=�'=|&]%��7#2R#O�� �%%Z ���e��|��ꇈ%�2t?^�����W*�ȧ���%��N�y�������G�O'LV�hـ3d�ö?�����y��B�+�
iC͋y:~Hۼ�2�:�)�qۯaێ|ɚx6J�ٝ��W9�p ܴ�gM�u�_�������x�zB�e�V����ng?�%��Ktz�/�V(m� �O�U93n�JܨϟX2��S���.25Zq���X��ĭ~��acO�c��_�DAnY�ÌtȹD%$x0�{�u@����2I�_���GͰ=L�������d�j����ef,�iW�%
$�X��){����+�3����V�+c�m˻K0�V!����p��233�^Ċ��K�=gd�]�3oJ_tW��)�dm���O�~�GZS?��OS ��7�s����uDb�@(Xo~��Heڞ� C�1��Ȏ���*+�i�"��~�l~Q.*��Uݚ�'���u�,r9���P�JmT�vn�j2Ӎt��(����2�Tn9l[.�!p�� 2�6,!U������=�����;޾P�
�%*����N0a�O�~C�c��wh�!�sD��L"1w���ֲ B��?/q�����\L��Lu�A~�1�B��O�t�u���I����e��JBK2�װ,GDș�m	���D[̉����:��Y!V���\-f�k���H��� ��|��]���U�� ��+[���^���հ8��]��W��kȧ�m"�͎kK���o;�n�V��hH ��w��܄z�$3]K:�1�h'C�w���»�}=��IpRQ�E+�>�GW
���:�D�{�,����~��r袇�/�����mLz��.M�@��ť1��N��QOdA��J��m}8�SJms�h�5�`����."����un��|�07 ��'��w�8𹟂a����߆� �"X�Xܚj��j���.�aXW�Mήul��֤	���?wc��Ż|i�X�FO�s` dL<ň,���nNu%�L6|�����7)-UFn))g�ύ��ZhMRP��l��o��x�s'�Nh�8B�#��]�����3��O�wݽ��~���7��AG�|��m��w��a�zq��f��潉�M���]DK��E@��&�J�������{pb�"i��7�p{U��E�ɨ3p��m6p�����vi�yS����z��OG�v���u��Y�3�[y�<�}0Ɓ_p�a�o��-���7G�T��9}~K��e"�����`�D
e�ʬ�$P�.n0���~m���2H��޷ ��^�,�����@>�[����M��U[�hπ��՚��o��ˌԕK��g>VJ�$L�c���l/��E�#�/�aŶ|QG8m�J(j�dbv[,ة�aXTo�||��t�錱ւ�[��k�j���xr���΂�WH�psf�0S�)>��&p7�No�o ��$:����ɵ+�d/�z�@h�����1Ansk�h�6o�n���
��١Ct�(����-3R�[=8	���G�!��-�y�?��8q,I�F��Xܕ�lH֚u	?cuD�v#���z/�z]V_����ٞ��u�7��t�;��m+aDE������.�F{�#��<ݲ���{戃`��z�91'$�0i|�z�[&dWW閒B�nn�#L�3���kI�E;�X�i����&�?��2���V$d_��P�J��(7�hF��<�EX-���mC�9�ݼ$��>�_۫�s�f��$(`TL-�5P��M:AR��y��_ײqmw�MojƑ{i#`�q�F�15�"S�G���c�~>��7-уq��*\k���᮷�G&c$$gɢ?2m����%@{�W&n�m(�:��+<�=�[�LQTU>J�����d"���~a훛S$ӣSc\��[�,���5��|e���}/w����8��r��#]����E��k��[�^sU ����c^q��*�3�	8��@��S��O������IV*}�-d3��+(��8yOC�3sؑ<�� ��z�QoH�3K{������K�n�wb�����؋�%s_h�F[T�Q>�� �Sh��.��,���Tl;��
l��r7�?�ͨ�!����TD˚ӝ��L���6�	C�3��/T�L�-�.X�P9C�:��{����͠�E#]��lVu�6��v3��6�wr�5�|�Ox­��L
��|����f[� ����E5ٟ�����UT�8RЃ�������}�o��@A�����P�v�$�f�v�Ba\?�@���ۙh�"���*¨��w݃}2����>�:֏�){,<�Qe��N@��Wxe�k�Ur�OL?�0�9^a��ߒrX�pvF��R��1�5�=��.�!y��p:��Qk�B�gg�N��bNNi���k���5�,����D կ����ǵ�����5@�>���+�G�2�����w�~GN�̦�4�'���H���h�4���� �?��>]JW
~��:�M�d���k7G�����K]	���@r�/�.;�U%�l��E�D�Q�"����sF�G�w����E�DŘ+\��`��+U�5I���V�Z�ޔ��[����$�z�W'-^�*d!O�/��tG�?G�=|�O�b��h�abZE@'�W?#cu�C.e�X�{��d4}6�e��	ow�1��!�7�%�IzҒ�2s������M%�|�?°`�HXO�K��4�c�`+E)y�sD�x7Yc�x]�#�E-8P=/��3~
�*T�+/(����!P'6�U#p��:��^������pL�z}�~J�-<]�p�(\O-�]9wt��{1�M����qnV�7����tt=�xc4#>d�-Cp+��NHV-�����8ի�Lvf:rP����u��4:]&y� tR_g���[��H����Oi��Ld�Q��5і�Bs�+�>�g�>I�����Zaoh������%�.?�
��E�c�A��]�xD��e��5]���/ σ�t9
C4Ρf�F�H�*��zr�jD��ZH�}7���a��7>�n�bvO��ko� ^��W/��w�-�0�̏m1��9=����a /�{�YI;3B�m�}<f:m�A���8vDrQ67��9=_��f��*�$o�:_wG�����\�r�<A�;��>c<�ܑ^�aCxAP��"����V��4�S6�݊-���������8M�t N�����^�No�=��:�(c  WgdaI ������ŵ)>&"~��g.� y���^@[��rp� *}�W��_:] �zQϕп��;�J����(�ڴ@�o[��g޹H�]�x�����"�M�D�ߒe,l�K^R�k�:S��t���8U��ˉAw�˛D)�z!�鯝A��*���tA�*΋�쮉�A�S�A��,kY�~.��?��0K���y�q8��CG�]C��/sA�f
t��s9	N��Ar��/ ���)x׺�j�Y�^3���Iר!�T�o1$0�ٚ���:251����x�IY�Ƣٹy�NȤ�B�����Eh�cT�N�D�8��׋��)9����$��=�(�J�5T�������,L��������P�(�(�P�t{��sn�L�iM���zז�zD�t>�� ��8�sͭ)����a ��R��޿L�蠢{6Y��%����a0%�H�W��K(�n�]���?2���i\g���w_�چ.�&���mI�Sf�W������\a�K����ɋ�9�)Z�	߲�b U�lo͌D�z���X��&�� ��޾���r2���+���wA7�NJ Mɐ��d-�R�Q�D����e2�A�e�}6��Z(w$���U�p�1��e�2s~nU(�X� �J5}1n$�
䷺��Gr���Ff��]\��Y�27�۞in���"D�k��X����Y���ݶ0�su��~Iԯ��D\O<�!�<[�nȂ<�Ҥ�SȖ��ڿ�%2�X��@*o��c��a{�l��SuOS�����_�ߒ�o�Tjߵ跏)�'�R-�����uؤ���Z�.��!�5�<�[��f4�
}q{��_�H�5z�*-��7����z�e7b��z�h\#ܴ!�%w�} �7T�M4��*GIU�%���?�=�R��g�'��n0-�kIf!ɴ<!IŋOҹ������R&Nmwgl�ԯ�Ǆ�؎�)YPA1r�L�Β$�[�pWz�ͳ�hm�	u�\yt�=�fd�
���=�)�߿A����ݽ�;���H�[�;P��xK,�y�_���r���fs��EVW)�.=�)B��0���+cA�e�Z�)�M4 ��F�oZjM�R��d�l����Y91x��
������Qc6h6��qd{3�b�J�d����TI�s1��&Z�Q����C�z��=�JEu��,тҝz��	����?,�{U!29���x,��4x��á�w6�,���k����[v�����*V.�!~MUu�<)�,|�AQ�m���c�-��7��~��I��Y֓�����$	6�4�7�7�G�$_0@�o����gT��Ah������k]'b�[nD�je�:�H���[��y�!K�Q�W�T;$�l��z����Fh��1J~?AD(]���B`��Y���y�wy�d����V��µ���{v�#�zڼ�:JC�҉HGC�B
c�x�DW	F�!�}�}P{�L?����S���൥����%���(V�k%�6�������!]Q���v�@���z-^-7f$P���G�6���%�P�o�G2"q�r۩�}�ӯ�K�S�'������K�h�u�4)����y���
R�F���c~�f�4h`�_�܉Ěa�~M�-�z���@�8��q2e�����V�Elj�"��u�a`������?/��~#���a��ei8,�bm��GW0��!�[�N����4��E�P6���q�v��|�?p<˃��t�k_�=��ף1�J�h�p{�(�%�/��/3�yBu�7XC�i(�R�����a��c��
�3"���I�pk��\:�G�����2,��Y�5x�%����X��d���s��ץ��Y���Ɓ_�ɉ������2ɝ&gE?�?ꦎrL�z8^)�����`41�M=P/�L*CE�5�u`!n�>.n��߀��R�ZY���WQ���tMݻE\umo��{�4aR~U)^��ZA1�?��\X�_;���g�e������L�
�����Y(��9v8�%>�.��r�ky\!W�$�Y����a��[�Yc�I��h?�����
X�������H��B,�
A��p�F��'�X~N2�Zhw%���0�	���asUiB@��Zկ䖩~���7��F�_
N��X���K���5%3�|���|�2�<rb�4P���;���-�+Jr����j�Y%�8����A�y�
��|Y���F��F0@�\>��T
�Ԁ�rjd�����0,>�>D�Az�GH�X�iT�e� U\�uI�*������WM~%J���7(�A-����N���c=VA#�?�J��2�G�Px��aR�w�^��FZ=�~���Q���;���k�[�.«x�v�F�؋���g�gA��s*�̊vGm<X�b=�2�.�C̤��t����mH�E����2�Ϡ��,���,tA��lB��h�)�5�Y�*��³�c$9��F~/������3{��:j��b-xt��*Cr���#�z��8�+��	kAe��_}�	��*���z�;3��k�sR�M;��E %��!o���iC��J{�}R_bkb�2"�~�Г��q����,�����:W�OkF����i�R�HJcv"� ��%����z�j�+
'���A�\����(���dE��S5q��gd�H�k�X#�c-��o%�<i�!�� ^)s�����>�Th������e�^3�`��c�b�k��8�M�guε��tre4��V�W���#u��S]	�`X<`�1�q���i��u��up�P�����ƻI����=��*��P޹N��{�1&�%w�� �����\���Z�3���z���%c"~�/Ŧ�~�JZs�dN˃8D�A��D�`K<E���{�E���0Q���/���V��y��8D;ۓ��#��AK|�k[�'�X����I��'�N<����/�k�ċ�R�7N��t~xUP����/�\�ğ�^'�ע=�s׿�w�B���F�*��=׫f��Ę��g��4N	5(N��=�6��	_i��c<\�������Y�|O�K߆������ߟ�~�}N�(�;v�2�seƷj�;�������&�B��ʔ!g��r�@,C���U�#C��I�M���e�C��UU��"����v�=�ePM����g�fsI9/��j�u ��T�����j�󔃩�-�*M*1EQ����d[1����I!z�Q��p�(�Â��)7�w"�On
�*R�z�1���ADj~i�V��zc�m��].`�O�%�c�4J/Ꮔ[���"���F�'얪[4ի�2���?2�Ŵ@y�yD��7eg�����C��b���_��Xt9z?GU�/,���k ��St�۴Ң�Q%7�Y�l�(d՛�D���0�7h�D	���0��[�G��Da�WCy[�o[Ў�Q�[Iݮ�+S~����}��6�0v�M�%�e�e��������ڙ�pw`��v��ܚ���=�5�A@�v����6�^ڏD�����UҼ>L,��es-���n�|�dm���ғ��Ϻm?�+'�	ܽ�(��HO� #��l�,B��g䞏ٙSS�䡍�:~��T�IA	�v.�2�qjl;��W/��C���73�3�+��j�i�}w�*�/G�F�>����\V�ca�[��4ɫy��YG��ƴ��`6E�\5����� �‡��\��&�������9g`a�VܔeǮ+�⊵�!p�֬G~���!4��}.���Қ����}���D�2fMd�͘*.�c��:ާagI<S�*���E��@z�|o�3����e����8�����a8�6����_N\�����Qh�����M+kt�n�53og�8{eaDB��X�Ńte�x4��ҏ�^`��1�������c`eo�t��Sg�cz(_ؔ�'K�eY�*�GU0�WY�(���5��h�b<�A��݉VK����jju�(���nS���?�Ẅ́�K�̢����l��b2=�H��.!�\�9nZF�`�KN�����X���<Zjp����1Gߛ�,�;;��
Z���FP�ѭ숭{*Vx�Ly�����H7�T} 0_h���N�K������av�?\��G�J��;�'~�c��x���R�Cuh���H�U6�}E�1u���~%�T���i�ZOUy/��(�P;�ۺ�%�v�T�9ɿ*����5'���/��%�W�!�ҥ�(j%�"�ֶB��e����P�uV�D�n�N����D�p���3Re�2��/�!��ft^k�=kS.38��V�P$�2����o}_,�0U"��Q����nd= VJ��I�>+�w��g�����L����!,٘����zu�J!O '�35]-<'���cw��S�|�=N��K�!�V1q�&iDc	'U�)�Y����1H�%<n���]ݻb���a��h��׋�.�t�����1F	���P%��ZD��A������ؤ��t�00˃��g�P�7�4<:j��k͔Ң3�WC;��`�ң�5�@ҍ��zkqo����L���ZtB�I=XMt_�r�L+��25P6A���^�p�i�t~�D�D-iw,��̝1��og,?OĖr�2);��J���,:1��si���V�4�0�b�{i�F.����+{�;*��.�3F��@��+��[F��=q'5���y�<vEI��$����r�d�`#��k������I�����G��{v��;�!���t	�2A�jݑ��W�����Z����}6�n���T>�)�`g?!<���@�����c0�3o�k]��ZpwP|�� ����T�y�N&�V�R�K��B�ce��ȯ-�3d���U��:�/l�O��ݜ��9<"�¬!#o�m�h���H��(J5O�C$�`}܃��u������,uu���e?k��%��Y��H��&H����T����b6cd��o|���[����� x㵨�rȰ�u���M���߲�N�l�.A��}a�Ukc�h�,��X��h�yA=h+~ĳ�Qi�F���Aa?e�8l<8�[���f��)5��S����B�0�I�NC���6&��3�@=;�H��6i��M�XbK���3�DF�U�}c��J5G
54}�b=�oi�ѼU�~!�0��.^i ����
 �>Ayn�����@FY'�(r X{��1�FJPO�{i�q+	����n�mѮ7��@4������}s��9̔�,�Td��Dz���@�)���T͋�h�խ�Ƣ�G�7u*z���cu�J9����E-�pO(Ac⩵��RWF6o��kSCĈ,[xy�rz~��C�C��$Y,ȍ���nR*�Q�mw���y�E��VēX�� R�7�r��3���C�c���-Π�lcP���a���!/��c�pՍz�f���-V@]��Auk
e�$�b����LU@1����RP0�����H\ΰ�#*|�u�y�D8g���\=�t���ڲ#�?+�ߜ�xCC�&�FT�k(By�:�̥Gh�p1��1K<+���6�`	[\�C&��3���I  �t�� AΎې�F�K%!�m#01��$F�-`�0Sf_R�C�8��K]Tb?��g�b�Mk��ށ��T�(Mbjks�l
$
6��K�
#ĭ�[y/�"0�sI�e�(Tg|�>��Y�f%���_��;�U܍
}�_U�VԗŌ[���H��YM�@Ed� ׹tl{����t��5����=�Yy�#�_Q ��~7��&����{�������J��[���n��gJU��,e �	�{�i���c��\W��ۘFP�� �o2��M�����K�����Q��z?==�1�y��ckt6V�ք5��y���6uI��L)g�h��|���D	.s��}޽'֬�7*zo�{���?3�y�(լ%�Eѷ�)?��D&6-�/���3�f����n�C����q���k�?�G��
���X�۰�r����CcuR��{�����8+ ���"���B��pB�},N����bb r��|���D2{��'R���hr�";�p
U�q��&�̸/�@f
׌aͤ�")�H�)��g�T���#ǎ.e���h� /D�ПvrQ^�ȿv��C��Q��y��Hd:k���<�T��J3)�xFxCḑ���HM��R�<J���c3�(g9#��tv+�2���ӜZ���a�y�܍?~N������_� *|�����	�X�������n�5]A�!1 Ɏ�\�@L�t��ꉵi�z۰��6�ͪn���Λ�N�[�g1���(K���C�v��
��BpF�2�DY p�Ԃ��n�}Ϳq�Ja�~�˵T�ÄԲ���9��Z;Y�o'��z�����>f�kI�E�nͳ�a�h��R��-�N4�?VX��.���t��Yࠁ���\�0[�aֱ!��~g<m<QHE)�6��ss�WV��fI�Ik���'�5��8�;��7T�2��(�;��FH�G*NS����Z�l2��N%��B#�r!�3�e�N�Dll4��2O��v}����̧��'\O#=� 3C�!�D�$I�H���
���CXx+�N��&���E�m	�H?��E�{':/CPv�￡K����9�w�I�,�V�EN� ��a� �/�]���W%�}`aQw��u���Xu�BMɝF{��5�}�Y��\�yZOޱ�<����h$=-Z�~�M{	x�U?ZΖ���� >u��������ǲ�!���ҿML�䓂!��G��;�o�ob��=l}��9m>wy�	��S�
&m�f��'=p��RT���6��5��Mz[�Qf!l�?5U���V�A�`/0����I�
�b��~���Ӏ�}����fn��� �4�{ ��+N��5���!�~y��T"�\|,�v��5-���8+�;�s��e�9o&�KjQ�f��j=#��z>�x8�F6
�l��~5���58����)]_N�;)����x(������� ��y�f\��1�"�h"�,�-���"߲ㅝ �����Kh!E��C4������)�qJn%������޸�~2F����� ��Zifr���12:k��l��Jp����<�6_EɀBT�4�q�LgJK4ON�,�䂺����6��y�jÆi��t�8�d��Ƀ2�i��}Z8G�Y`�cOT�I�аRSl���.&��N�+�M�o�����t�90��<�j�,u�7�%����̽�c��.��֏U�<�w��+_z�ߊ#�lk�)>,�&/�"�E:[x� �Ym:?N��"fD;�����,!O���+��&b�g|�+���a���?��]��	�|;?4���/o_�Wx�IzW�1g�(���k}��Y���M�M(�N��3t��ī�v��x(���F�VRk�v��ʰ5+t �������f���g�g55E�!�|*�A���|D�0���5�9I`��x���	z�ތ�C�N�+~���N����.N~�/�6��)GBZ	DV�><y��x�� mV�3w�	����ti���r��́R���@��s�-��I��P��tr�*��X�� �D�*.��AVU��Zy���4L:���0���O_�P�閾���@Y������1d$ʉ$<v�Y�@%���cAOI��o�+�-
��9�0���X�؏�2/�̍���kJ�Md7�������>���j�z?���kE��ǫ|��*���q ���0W1�0��	����=F9c�����U�Ď���3�u�u7>�X��K
��t�ӝ���=LM�$y��ԿƟ�f[qrY��hUQv[J!鹿_+={4�O�\?�T�ĭ}Ϭh�<[�>�3��O� ��8�W����+��D�S-�I>�E��GQ�>��ӏm�� �@��rC��7�ڶGh#DĪ�H@�����;���g��o8e47xe�I�8g�Z?��Q��cz�1�HHU<@���mE��v�q�۬s�i¦�=���x�vy݃0E:Z���6}�~�Cx.��6���:C�R���89hs�æk�(j�����r�eF���:3^W�x���P�x6�?S�m���v��&�1����<� %`Q0zLE띙��]qdl�i���%%ۄT7�{�)'�MIkl*�����I��	�-w�~�n5���м8���J�S���l7��Ū�ׅ�f��8T(myX�W_�N�l.��·<�[�|�j�ka���c��c���e��yZ0�W���)���SOY���p�k�a.�En��:Q֔n�g��;
�a�`��D�?�&C�w�������VJ�B��3yf��GGk
A z=��+�k�i
��)�:�p4��l�5����t����!v���r�����[Z�+������X^��a�^��cpb�Z#hU�S:3�=d�$����h�CG�S��}�k,��?�a%X9���T���C�n	�-%�b?1(l���t��	#�:|{���4u�(��Kf���N�JI&S�
�(`�{+�zR�-��t夼׌-��L�ٿ�����>i��-��"���l�-�U�L����� xƲ��W��b`��q<4��׮�2�n[��&t3�]� ��l�+�r�qN\�z�7Z�H�E9�@�)Q0�}�,s��H������՗�hY8U'i �O_c�vL��Րy���Y��9��&F��Y�\q5���48�pQ:3y^�g��_�8vES.�w��-7�_�"fϳ�m�O�+]��"E�J��$k�sw B�yPć�)MbhI/�a��P���Vǩ��@�<�Ѱ�K���K����y5_�����m��ǎW�P�-z��<��>m���H
�c��c�c��{£�� �k%�����2�ml�CSm������&Q�V
ue���g��C����8���6���@]�����3T2���g:.#�¥�(.0��+�����-�E/���:�� }N�|.�����\ _��;�b�޲ �A�W�+�����8��,�kXv0�+�'c���E-��� 3H�a��g���T� Ͼ?_n�w�G%!�c����yq�^�aq��9�H�#��Ζԁ�	F4g+lI���2�)�j�+G�eA�=}��6�*s_��`��Z�ϟS7h� �zU��6��|H��X������#jb��6)�8]c�T��3�O�����V�_Yᔫ�o[���f_�c�
�����9't0��.����,��������0���>��JT�*���fo�ľ���_ʻ��������@����Uf�����8ƽ�^0�v�e?��a�$ry��!N���A%T		J���1HI����{dY�,�Jy��/�PL��������+__vB�]^��/�qUfe�&k���E�%���D���p��}��k�{[ �ɝ�>�S�k��N�:���}�X�`�p��@M47+�6�M�HJ}G@l�b�;i�� �O:����}qض���.��bF�z�~��i��MsW�
ᣚ�z/��Wy�#B��d�3���P�{°�F�Ŀ)��mb�����MFY��a����y�@�u�eJ�iDl�H��#�';��H ��]��G�vr�:m&ysb$s�_n��V�X-�].>��ǒM}�Jp3>�_�Z1��Va݆���r�.��.Lſ�iuTsgd��
GP��gꍮrb������?l����ya�nb��!���o��T޾6~E"(��In)!(G�6X�{��,�Wc����z!� [xe+xvˀ���(0*:l���ւA���(:�{�C���3�4s�Aօ��T����Ko��Ѿhڷ R^R-����F=��p�	��U��a�_{��l�bw�N�f`V��1H|� ��͸���gr�cȨ��a Gcm:����Z��6hќ�܄�8��e�?�f;��c�q;7�&��K�Zbr~�u,��ǹ_jژ��b�A4�W�
�����I���j�K�\�A7��e��]X�H9N��/Z~hŅ�	����d��,W�P����������s��&Q��.�b3]d�:�2��d�;�����?���©�_ఱqmb�mfWy,��\$�;��p���t6{�=[�$kP�]&��*��
o	c�;_����Gs�ҍ��s�n�	�B�y'�f��ߞ_	AL ���\�ZS�W�G�k9l�V�i�Gu�%0k��׬R����eÑ���璕K�þ��v�Q]s��d��_ Ex�|�;�z�*M������w���{�(���qk#c���#F �8 f*-7�J��ݾ�铊[_b��_��Ð[QTŐwF�m�p�w}� ���u�fR���n��˲���f�?o�r`G��TBV��Q����˘���֎'�@�:�q�k�1[x�^�}�T���v���+UΟ��
&�U�Fc�� 67��y�TH�� �ϫP�4��^�	��#���S��t��T�Xw[wԜU� �U%BE����2�m�seM�7�~�����%-l��T��6������P(Q��GW��.��d���������}�D����[���|n,
�pR����]aߠ�]Y�Q�#�?xwO+����F|ε'�d��*ߑɕ�O$��`(U����0(�&�*&������P��z�������08�I�<�^rcss5�[�`ў�~-�T91�?s�q�5�N�I��'���z3��T�S䥤W�O�@���:'�jg�G�b�g<M>g(
7�*�)��V�E�5Dz��9v��/�g�T�2'�f��b�]���KѬ�'����ד0�}�� W�e�@L��͚����:`.@�<�J�M�ho��E�,3-�����"O���h��@ }�K��2��[��ٞ/����rK0N�#�[�*�r�7�~�07�!\l���!lcV�7j[8�6@��-��Ｑr���t,߼���%�8*�( �T򛘪DiB��:����;���5�ʀ�{K�uU��8�a�� �������%��l����\�i��!�)�oY�_h��z��eJLXeM��������s���u�A����VF�F�UNO��!�	�EV��Ȱ�@��AyE������������M՝2�`$I"�Re��,�$�a_�,:�xf��ʞ9����LK]f
����~,���Z�q����߽~�j'�=fT07H#@D��d�$���|�C��������ai��,�����������љ�ش�2��Ҁ>|��1���"L (�3��F�|q��A��s����dT>�����u�����{��D�8ţhذ~�T�QPB';uu]�*ƪ+VÁ%�i~IK�/d�����LZ�Y�X�حI�K�ڌ+��k�f�e�sޛ��I���݀�t��A�v.Ђ���0 #O�J��6*�d�ēMd�S"O�������=5D�e3g�r\]��H<W�qϾb�j�2,��|Ⱦ~�'���as��S ������N݄�}�c������j����n���f��2��[�JR���Y^�壣�e܅�hL9��~�,y#��〉O�}Fx��t�dА%��Ż-L]5�B�p>; �P�h�}�: ��ɜ�Q��6*`m8��&|Ȱ�`N��	�~ąP�F�������ʏ�|�!���⢆�F��Ve"��^7{1���r�����x��G�|��UAPM�%��@C��BֹPRC�V����Tݯ�O~i�d�*��U��h�I����""?B�o�ܺs
�d�X�%��y"����'�r��ok�Fj���ue�P�"�y-q�����y�㫉Ɯ�=�.(��������kxLA��ZvZ���B������6��6�?��71h��@0��&A��J�]"���������'����؅�(|"��Y2��}۸�>^�
#�����]�c�͌��.���$�'QQ��7@s/F�?�����t�D)��O�� p���޲Yn�l��7�H�� �I�uޱ��z��\�c	�vt�s�E�+�7vt��;V�Ls��o:�#�+��L+=�/A?':�i�E�@{�,�I5ǯ"2�z����:�^K*��Gf>8��_�-�B���9�W�weR6�`�W���a���\�����}�؅	�Qv'��5^&cէk �I"֯ᅔk��Eh!��诱C� ���si'9sb���a[x�C,MI�5S���&��r��y��զ�z=Pϕ �V�/�+KjD��M^���z}���AvE�.�	�[�'f�J��h�q��<6�)/��A�H�Cs��~�U����)�p��oeۮy/� K;o���L�d��I��<�r}f���H3���C��-�Yw�;�r�8l��f�Y�,Ǟ3GM�y����45'G��>�������B��q��#d��6ن��f���6jYYgVm�2����o�Y]�I$���Ksd��@�-�3(�o������f������|UD�1���7@�$�ۤ��p��4i�+-}V���$�o���UnK@�{�S�W�O_+�RE��yP�bbua�gS��z�M��D��D�t  ҥ�ۻ�.A
J�:XN1��pc�˝��p���P=5VП��!��=��/Ƚ3�q���tH�&�\f�f�[ݮ1����Y�x]g7�z
