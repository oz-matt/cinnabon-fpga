-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
S6N0rFGn7b8SM4poYXHQvzRxbf8gmNkTgaFSShWSZ7pgkwPziSZWxThHG6Bf3nqU+mKUEcc8mebD
dgw3yxalAqeD7kByzcBVBtEuxc3j23LAZNNFB4RukEm1H5nP0MUSopOEETEmDa+R6Lxl7plfnP+s
dfaTi8/7cbkDYuGYstzzyDlK0VcSCuVRjVnm59ZIH1JwXC4aPdg2YeQE/DzP3SQYg+0viqBLwcee
ODRAxNo65D/d9TT2/Jykrsc4W0J1Ymvu1jz8BniwLxokYXtZG0OMQl4e28tCAbjZXG5g24LTCzlX
ETn8XHfhbmeIo0m7USwYEh7p1TSDM/ePdYC6Fw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4256)
`protect data_block
mRLk+OSfITcNOIoyAwAzw8A8D7/CIMuaMNRTrsj1UpDhWE8dObUc14Jg+gijyGwbI1LxqQs9SJtA
qdWOqsK172O1tlMbkHlpOzk4xDugplANe+zJrqfxrXGmm0OX4W5tMTZdSDL7CWJ3Ep2Fu0/w1j+S
ZRwWHV0BkhH4JdQriq8S0u4U/ok/ecBQi9+feD28e8IVfIKd6LqJWoz5dU/mXKIu5ZQSVYFq9kyZ
ZdLRlnp3UUL72EjR76OEdb8c0NNeUhMRYpUpkzKtiwN9Xs2tQ4VjScx/QoPc94cg0tFRUVgTKDVp
IZ0Nfi4VPfV4sAb25kOPuWKAcUuJ61XU9mAp+9HsxOzLGSD6VtjdfdR2kPEjKFjMtmjs69NksmA8
XRgFZ+xTMX0xO5b2VMPem/xphWVDspQlZ82UKjkiaPRgaKisr+/BdXzKBS0JinSJeRRCbCtChVRn
Z2929R4iP1ne9bN8lpyvPcOgyXJ+NdEtpnm6s4lwmWpVgGmDnE4pwAPLYVdFQnFeopS71tThD2nJ
M1AdCeJPolH3m7qYJqVccwjYk26QbgozHwi0xlrj6awyS6Ke7zepf96uM2cG7Lkx9WucfHTe9Ogs
bP5cFyhoqiABcR7aem0pHUlxHRnv2mYi3cHrOcGev8JDN0+vllYC3SPoainCRCtS2o9F7xqH4CuY
cjCwgOpJdLVMCGVFBlZvku8ssVs3eCx0hqiAqFxz7xmF5xKcz3aZJFD4R5D9ROrYaHMkfXVqFnZ3
epnkUbwzovI8NjXItAw9IpcUkM4vE85cSyi033aYxoGty2+bLam0a7EysNK0vJ97ApQHYP8iHaMS
QoCH+dc1aGQmDb3t0RcDwLRKjjLYO+bfcy6/48NQeJaOJyhdV7usbP8GwaXhO4+pODABDHRPxOh+
gaeY10M54Nm/Wp3N99pgv4Bswlj1AoGR0IpbBpkSajVviFbygq1D5SvyQzTiU8xn0TCZ7iouNg0a
kmyLj4pJcKpRzsVp72e4sLwBU1SBliiTz5WDYtcrFHamUcndzS0vWXBWab4iBPVZGbrn0GGpeGmi
NF+8H116CIS/LfrIEhQC87iGECq51aA0TjsvShyqDpqDA/b+zWGM+sJ6S44y9qexBztHMW5soLl9
E1uQlJRRjyr8zZRMJkesVkPNjEnPPTb8DezUu0lp3Cu2KvLiiw0MOPJ5M2WKV7LQCH9OxGfwVGwN
79mmPZWTFwF4UUwMbqilaKHrhCvIKrahSHvOrZzdM1YmbAFrhc4j0mDni1yX0k/p3z+6HLd9iGJE
/hdUK0U4O63JOIGcyLxjtp7plyr3j30VckN/ZvErOvyEgV1/BgwlPftOWA9J320SujO8zA1ZIlpn
7e4N5kDwcV8Fy8BJGzgzIe9MlnPg/VGjvR+dEEk0Q/CFDeVurnUkr1wvrNxJcDUkBEvTvHr0pHfZ
/PUfnUAnvkQxAn0Gw+ZJsXV4woyj7VeMCiDx0VWwzjyKlgfcoHTZQpD0dct+WhLlWv0ICYK5dtKC
YqioooxUjIkSXyrKsn0Muf5Iw9Aiv9yQdD2Wx1hafXfB6n2Q9fuo842wu2T9c1fyR+KWnYnoAta6
yIou9i1dXOTccO1/EreU5OtO3YC2G5ainKAf16QG/ovfeZWQYTQXzRwB0rl1qbLIJwuMVGmz/D0j
xDWBL91+lomtAFO/qftov4UrbkrDPIKlbwTjFPToHF8X1l2BLjF4OpOKakC9oUVvpXMczVff9of0
vSls9zAYb36WEdYClVMeF5q1DLlgM3gdpnvENphGokWbOVWxkWM8XBryte8PXAbctvXfptK3zVk3
vWyrBPvNTTJCbkUdiJTbvaeU9SDl6Mco5KKQi0/F4iW/R6TuIFmtGs2Dq0R/8QAjwFLdfC7W28+X
GgB9VJS/DHqpOck22QcJJrC6JnlLDkXy6qfnyjoWvLFI8YbdfH1eN3TE/zyBEuAwrV/UqOibW1fp
3KrZzSt3jFN8rYsKy/KXBk6ztX7NytTWzwkh6FAAWtE2woQBlf84BmxdFHMUBcRI9ZsosHEC07yj
ZNmNb3eK7bcyX2ab5CRXzADxfwgrCjyxRQraG0loWiLtVVYiD3s1LzGI9m9+4MXGYKHWgccpw+wT
J9U3E3nJjSlZHw9YyVQu2GpYmb9H0iovWpmLkDWYH5E4wwyVd2ylvEaCMyejYzHWiUQZ7eu3QWyV
bAa5Ah0a7wT36GTh2ykiQRDw9YX3luMgoEFVLr1YU/nqFpVUOEzB+dJPHLQeUMUtcfeKnv39lidC
+Jkt8h4YQGUjFkJHOlAFOAfA20fmebGsPqtksZkmyzva6Ad9K63XsrHvv6Xx1yCrUhC95CBx320b
xEl18n5ToTuo+QxyQ8QmoCXO32EzjoHTV2AATd4GxAYB3TUoFHK6vu5qDXrb89za4gvUNUpK+1Fm
5YsWxQ6cQ36GVlleLTQf9nmyROVygPQz6TJoM3KL9N2mFrdrVWpsdbOSfrLUks5rt/+i8Zxc1Dmi
/+Fdo5SEkY0S+e7+EElAP0oMJy/QvEHWkYynrDGqhsa1x96nQ1Tyomr8SBnpOts57tpzodD3rVyG
HNUXKFLYcmIuATXqghCHggtXpRg6CHYlVxgeDRE8F1etrMouf6jMlBvFQSVpLw9uPtDTT6wKBruZ
JbwXs2/Kn38ycyW2doaQCxMEX7k5+l7XAPWPWyjwGpNrCqr4+EJINdqTrIG6NkkSiZf6YwizwWVg
wg5LCPP2ZyBaCJa3SjsBU0TxGHtA3cM3LKjQBaix4JbqXXdHtrwX5OEFBOn0FwEewyDwRoxMcbI/
qEnIhPQnYHNBz2PSQVyfFpd5NMnRhAbyI6kjAr96VDQNvKhjBdfCUCMPiqpoMuZDuBK1TBetPKPr
+xcrjqFsB+5opUf/sRxlHJqydcCtRmzEFd5xk2you3jqsBCli7UsIWxEME2dlkERZNCvxBjdPRTZ
PdqPe50oa3EvWUWalveTgRx7PFDByJMDS6RdrbHBEnlt21lSAqaqWrWmiG+B00Z07RiTEYPoPrif
9QotsJoWQzXzhYGPOodxqkYLtP4VJPK5NQcs+3ZqpZcgn/hxz7znYUsGAk7gmK2X9D59iSvueyk2
qR4aubXyDcifNyDQXxwlpDNUMWCTWipQHqWB9ohCOgYxuBUDx6ntoa0tNedmKjpK/CJ7l7QtD3Xf
cBfQ2fbOf8skLgO/yIMnByyOLM7GHrOLgohnbGbMzIUBUFGvh+t/PYbyEgINld87kPc/L2LVdQTz
DKDiSA+uXw1bqw85PL9GB6x8qy6fOYC2IAw2Ec5Fw7/SuE0AOR0EYVosSi7l18G0z0THdXwfkATo
QDY2ORi822TAp83NkusdQqPrx9+b0PTgOdSd1H5n6vrnJ3XGqKkgMRS+QT5vmFhEKr1iWpiTr84n
jfrPSSC9HrNz+iEpfizVe0Puy8ayJuIda9dkbSEH3mAnltxiOeVd2cCTBe0I5vmqX95OObuklbN6
J7EPqpbpuQIjceetbgCxQYeQx4/saUYpDPQaSfdOjhF8kv9zFveQJytzGW7K+Q/pyIxF9Bo2q0Pt
QaGU4H8ALkbaBCr2lfiBnxWeLyZnorFpevyPjbwO/YhDWpzUxxiQdOiVniT/sc1bBkY9MJRPaKV0
8utVcTQWyE71Ac79/6gzmbuezf3NFDQaSnohMYKuNZX3bpqFF+mmslfCrEYmtseMJJ+hTRfwkV4P
HsUNGv9XaZbz4x8MFhu991Uep6tfjO9iW0hp4UvSt8g7WE5naYk2d93TUfW7C4yG7SBLr31nk6pD
wZMhMUempgucPq8mWSPwGSH8xATI5V6XdXM7eOXNoWvV/0oNjVn6XfHEganf9x8z4NhxqJJ6VrFr
PKGzyEy/rOd+ZGBj5L83t6vfMCPITB7VZw2WL/rW5onvAKB1/3MMYV0lIpHMnfYElm1DFvoocZJF
EXPRgLmsdO9uYf8/DfyuOM2gN/bewfq4QmCBACzxCJcvkkAxea37gmOw5h1f3fOeD6zVASylaVpZ
4xYc3kOnDHOsRRhoUgEFBosL8vy33TYnN1V3AcfIjajjwpLTtAriYgMP5NCGOtPRFUH30c5YQbP9
QZax2k8g//MrsEWJ6mL5Zjk/SXPCwjNeBe9V8nUwZ3gol/OdUP784Y5LC8iccKbBbDHW8zLZPRBT
aS1Eqpm6WloCDOtyf61ZSacsIoW37GINm7gjOKWCzCWpGQ9mrMRyUUeQSK12T47b1lowcA6JpbzX
UVt1DJN25AEIvB8cv0wFUfVNLRVHV/Ve/Ky+9GDnToOVMLAjgvIygCBljGFc0/qs5gP9ciDUFRs6
z5GfsMeX9OBcwUtYCfmZXprJY2uQTqEoUCvKciIUFRh7w7y2I5dDBZNti9XkKpiEoPltmZ5Mhih5
lC7rqWNsQhLkVZUoC48NJjW+S4pJLhfjxEn3nBgjm1uLCSda5DQtraqSXL4+p1AurnA/FICqgte4
2fwkPnacYrzxlFLi2QpvwF/I8kD9EjkwMsUPjKArHLnSWgbpjTJM2OseCv6I3KHku7fPKUPCkJcL
nXuAXAOU2H4kk4EqlfNmKQ6F+NFSluLFzwVpWWdWCiPWBABk9PL8Jvs4MOltFVcdUxGNlqBC245g
BW52lmH5+tSMUnTPoalrsholmM7kZm+ghaKInQXD5FxFRLu6uOegOTTYx/s1mIsXpS8R1f8cZe0I
3s+ckVezmh7BGcYXGFM6+AfEyPBf0Oeaj/t2HzMSg+4ysqL2pHDbTfEEwFxUwXii0L3zmEBSbzio
853L6QKifvV8Fmom90VAJM+YzsQU1SFbseSRCviY81inrESZCucEQwYCmaqZm7scVnQaoKlPxIyO
FHWJM5XBpvdOBftOkthLLBWzSUZLCz/nLO2ajE+VRGEgNltfUGXlDESQJmTC0zbpll8emLznhSoI
oGTSopTGHXrqhjpXxRHKK8F6EXMDIbgc/0/e4C7VWI5HKjWE7UwxmEGvgfxcMh3hBTYZ/YLgs/0y
TjzNswOc7a+vDmAoJHVt40kGfSFu0McI0J7pgQREfn3e92PRi3ESC1wJfdnZdaKX+JwXnfWjcibi
79pYfdi2BfDNTF0eUgGIwVaHNSnv2yP6cabW3Mbiaz+Mm9lV4D7ajThj9f6HACxaGOmghW7CVDDi
kg9EiPdbTQ7pzX68v03zc8B7pIXg0mEkuviEo95IAZgQ/CaA351OuHdcej/00BkUfpCktMbDEVKe
A36VWE4CBekZCXzHhV7RTr97u9ZpPCac/ceoti/s1mpAPe9lf6t+cMFBXEDkRGyTie1dqIKqfjcK
+BL9VdU8xfjQVL6xMzgoWcQC3M1w7ker9+TfCEWxcB2HqP7FfMEshyOBPtw0GfcvrsZ7ed4mIVf5
3wsMfEvrAqQkjyT6qrIQU+7hTWUhMAT0K2YHLnFt4sBVPHlIZZVhsUa89od2Tv2pPfmDantX9Yog
P/wDUcIPOil/90RGkM/VQqO2i2qZga2NIaLKHAEQNH50y7sHdGOIAAbWvZFRitMt3ousf3hquJjq
z1S1bMByrnxy0IKI/tO6YMVqjmr6xjydSi5sYEP+pFHwdxGL8mX/qnamt5qishINdMFN32hBwk2/
5NFPanymKqFYqd9Qp9nx0273DRSZzb9kU+SEs37wbJ1Pzjs+PHQ=
`protect end_protected
