-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sLjR0t+GUhooVsegAK0KPuoEvPnuLN0Mty/Yw5Fb1Nsw/d2bimqDCuSCc00wzSaZh4KQJdy/zh50
+Q3Oi3/zjbIvAtOuJbZuvirpQln6MO9CoZlhpXwNBv8WT9kBFMUulGMLsKGRoRr6lGQ8BDhbSh15
gCRUUCicoP8G3MhdCIDxrSRT4FRW6MP8L03XBmUnGxy5a9rMgz8Wxa8Ga+ikYKN3btNwyQ3tUGw7
ZuhKY5lLWNCw7Xq9KyTT42PM0EWvg2JTVhArG9zI38E8ZtlyBDTdmY5gGyvLLeR8BUrLfoY/MMlQ
gTzVgLtB+vSsnLrrjssKrvZcrVmjnw/o4glOgA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6144)
`protect data_block
9r4MXHCbE3vYgjOKKY0GB75/nYIzgb1GGY1zmCL4vpXxJfX+LTgsZCpqWCVXvpqr8mrKg2R83aks
BKUqGapr25DrZpgvLxd+vtw1sRFe2NKjBWw6WFqd2D75HWz7Nz+NGASlc4/ys/3ceGWJ4wJYrstQ
YKfj/q4c0jqq49x+okzMkaVTDkKdA8Hm29Vnojk0LUDyCVxnc33HSYSYlIb6OG9W1V/G9uE0GEOh
tM8hMPavljmdBH1KCQgzHTKQOvZBlNYsBoKTK1emznzg+UyjS4bKjLSglHrmt5WVZoSvtS8u/+aa
2Xe560uMrg7W+SFMcTiEuV5UX+cBGeQgWbz/Eq1Uht18ArP45FFmDvpzGiaRNocoAvowtIFOwiDA
lfM+6KPYy6JM/jyG2oz6uQDFq9L3t8SFQLetBu3uyEfIO3ZSGlajkuYA5Bnj/X1hvI2kKVLSwFTO
Iot8V5xvN9me6Sh/cuPDAMTF8YDj2LVc5N/hUBGtUZUCyxFYiZ2w1uxc9g1jGA0MzrSHQm/mmVBK
cwRb9zGvKBpBUe8YX/xoBg0aEsaYIBGR7JuzwAUiQcaLZf/c6jPIxoX8fH3GrIfN82c2/oMFXt7Y
6JRpPa/dDrlhbtKQcATIEb0ocioZ7rszynz6XYvcG1GoWfQ2aO30JhKFm2uKA/6nol3VA24JAnYP
J94wiGhiOegMfnJIIs57ZGRQ7Q/eHrY33QvAn+2gdeaDIbqK3fV472bf5Xub7fiFk2uX462FTPPN
/8TjEHaq5pgzcL8z3I4HjkkYG5SQUQ0tW4PZTkuba6dZJ9Kai/CYDgz04KrOyN8LbyO6QrrS0NQ/
ZL5vlEl6V2ODcGbNZuhPXwDza7RkydDONYIQ1uPe2z6e5nF8FP+D9tDTZM6l7j0zo6MPaql+l0jm
QoIvocRi2KXfqcJt9btf6wI3TLPeU5J/H3fhI5KxgdCcEQFWYI37ZJMM1zyLoyH4MQ4EEn2S16Ls
BkjmrZ450dfempN3DHmlQMWyJ4m+L2RUUdIQsbn+Z9QB6xWkV0UkqohsoNKIbrAdKzRx8PHrgFW1
XDsO5lyeBR1+vCNDjFGOcgGBa818XN7PG5WS+mtuzuU55XCbYW93J5k12d7MyBAOoUc8rLKqjDOI
ItnUOEdzzGN8/Y1CL75dHWEtGCGwN+DS6RW0YiSlfxzazwQuDhsAmV/W4XFMerh9/MO73sw2Tr3U
MrCsb1DTlqFOlsuaTqAU+v0Oyuy2o4pT+EswXys8qkb78BuAlI2JYrx/s9sztC001Kzu2X5Peow0
umHUad3rGqdF0W3x/4A384X+HjEw4m99yRrqH5Dbdh2TBN4tLg3SyW6I2UsS82rWr/L9ZhDHmpZg
ebweuoXJT31YxzQn0Bfk2GtT6HvjORQmCEU9gWGinj4vd7AolQqMEPqaRHQIeK+cPan6R/3SvqhK
tA9GkA660bNtCLgdaGpEXlLYGnGzkDpmFQ0wr+v6BWaIb40lpzjjC+A14fh2GOiJZIRCX/xjEJrj
bHNAtjLYIW42k0L0k9N+i+Hb6fV2LE8A43lAhJUSIJ1twZgy7E7+S4M52iUTrYukCiNM1/8a4dR4
rBoaG/O8+h6Q7jy1E5Bl36HeIDU0AYglj8rmiMNUIBlxwdSAyJX+U+1jlJbLLcf8dnwNaUjsLkIH
qJqcUNXtHakqpBslUMZHfOx9XbaHrVE1O8lq04G038DXZadAlsc2sKXkcRMSfhhotrq3bP8MI/Qx
2FQVKs4HziX704GU0Zvf7FazTQLdxRjaY/RbCnM/jpkIEk6zQ1qbbXGENKPJwf/U6indISpDh/KS
Hn6eR45bARP68hTm9zQUVL/SOyhnIWaYMTAiarrcP3l6Sv1j3IEuC5LOeOL4c7QlLBLXttPZZmh4
/9n7G7pCgUE2hyNj/5ltCgP/SwYN9Imh9YfCjOJ8FZmD9DdU2Lnmns8ld+xd4RbVGvxpv45wSvEj
DV1LIjqqIiAUWhpDWOHwwfmDzlq9CKA675w3L3/Uml5UNMCaj5UxrP8jv33jy9lXwt5aWIkFvojd
Kqe37OqdJfi/4/wZcSioy92YYPbVlcq/7O6YhinoUbPEWiozkL82KaLMPe+OKSyrm2FvJOOIMzvP
uEVJ8aQCZpvoO4YiUrcCLmnBsYx7m6/oYA3hsqFic0tTGhIfBl7W17JdC8UGPES373t7gKg7Fdm0
SMFkYf6kjznK6PA117jyqxbwdj1wVrNAWK1JWFESAfxT6xhTXOzZ+BdrBYTOrQoNZAogGqWdzKsw
R0Lk2I1WzvgjXf61n3hMPgd4QjMyEzU4pbIWdF65lWX+QAeQSplTr2WQ9la3CIg+W5xzFBQGup0o
MRl4sgGLT+mXdYIpBOWwwKpT+SXES/bOSTqiPTPL5KUcb5XDSkCGDbfbR8qYvivSBHfOPKy680TX
k0CbUP3aktE/TV21dE8q/LirQJwOqZxeZn8sbYwYJVOYf/FBZpuY61wBmJlu9MEqTx1nICnAa/0X
UruWjCtf7pJ60+7sQ9aVcgFWVCCuFGqjBr94Z8yafYuXD5swMLer1zORN6/c+ub998tmf12EwkL0
CjVD0G7fe8ibjL2YkCUymr5z9tjMEItMMiwm3tDxgkfLo88+cqSJivm555r9S3JAmj1EVZ4YUfmZ
aYlgdBE4jDub2FNzt2wYyqhg6V5YKGm0u47jvBdxwDJfMF0MPsRnNql1rAFd1dJUzqyFAbpWWQng
RkuuzEEoubHnETXJsOP7bneJf/YcCsZl8V552bLY52bQzcZYtnpP334C95wXrOTK4iJUt0XZyoip
dK4vqHaBAjI6SKLfChz1UT5YqOwUCjnJqgWOCBwLoVvk3Y49LSu7Tx6IBilxYmRNZzDYr7rUb1BY
dm3VnzZ1lxViWAJxSudEAyFF5ia9v6TZL666f3/H8W7VjgAigKFyZvDiDkMjAXgBr3b7pL+mYcB5
Mta/yCvPK0bmg05Z0XnXUIgYKr7knUCOGIJMZtdcR5qWwkYUg9NNM0L6lgJ0mUb+TjT7tua6n0Ye
iNKRPdpm7+mxBhipal9TMu8mROW2MLUR9eT5ahL5oEloWqd/XDT5KuYC0YSnNW9n4vO19hluem5B
BJUvdA1PFNKy5bI+V8bVybMQIb7fzfk87zGqlP7tnYnAz0lnQMM6DBN4p0yRr780IAwAPBU/u+/i
5zVD1wDRu3VuxItfxhzlgWv9GwH/vfhKu6UHtAQ8uzZLyc7o9dMmPSWccaGdvNfhhbl64RNIuMmH
6P+dgQZmZ+2q2s58aM7kiPFsR9QewBuIt1kiNN3kSR7TjSJhbra5A7mokQnNNoVYWTKPpYG3sKCv
FvVJGm3HT6r/QmvHSGnw0xQXU7f5lAITTlVm3XV2G+GXPEP5ZVWSw2dbW2l5QtxEZQp3dSES5X//
bK5VgvZq09Hl38Zn1BOCD8qogxqCy5VL+fyw/7tOwTCJKpubLP6MtttVAUl3/HWlxu5Si/aB531F
4T8YCWPprh1IOeWcZgCmeuNNaO51AkPxAxE7ehvkl1DfG7+tZKJqixm/rpkwygNV4+N3Z+kN2HWW
MnOs6odI4b4o0dIxDdlZ/DSzPWmCToC09wy8y7x9FhcC9oiVmCZY70v9EIanC5JQdcKdKlzH5sbg
S/XeO0kFeJ04KtXVVCoIytFN5IE4GPsMzz9WejwQqTZ9N2fffGxZyJnTuCCSK4doRkX+n7ntDnFs
1r2FrWARGZ4dFyDYspiVpUCKLkMMdKw9imaAQTvQp8biXs2hPeg6LLr2RIam3xFdMmhqidYrH9Tr
pRoVNvkDIDVkxwQIPd0guyYRiZMjhuffX6flXtavn9LpQe7DscMO9XP205eNpZY26dl2oNwAyJJ/
I4upn4htGmPHf2OxK7vmMcvSc+m0NSc5gNFc3TaVWAaDk7OeE/Dlz5vkF8n0ECVbRV6zl5l+rxZ9
6FyB/9HExcQt08hpnTOwWzIawLjynzrt+L9mrvGWPJKGwbZZ70YUl1WWBx15I21Lyn3TGGm9HA7W
kfs5PvIH3WmEWM9Xu1wItfHGfzBHi7Cf7kTrILbeegWbUqE9Aa6jTlqYjDTQ/TxZZ+Vjn52K56hq
wfil6lU1VJWBQZE/OeWPbHXUlgx8Zp+muO7yh7FkXObZ5DGCVStj83ScWVs9g4aQwIkwyrXFMfQV
rZcdOWP1auEO2fQpBxkDsXBpVbDMZpNxhLmXAuhdjNTzdIE/rXRdwqsekhHwS16rcD666e8GMaLt
fy6Keuf2Gyc5Gc9PjblBZEsZ8IrgvrQYItqDnDtlQEopsjJ2ovEWc5kSPJVBaehShDZS7vZRPtZc
w5UjkPCxMYDLZ2bZbGtnCEjMbscss+Uz71aqDvXqQw1RyqOEmGr3vGWAlFbxc9oIaIb6BTOuO2gj
ww9GPAtUoCXGY8ahzhcIUhAW/L44zyMRn2xpF8imIKZbNkn57robjo7GPQLeWkaoail2Jn/XHjgD
wxSrGyaRDJ75cuVtXTovvNenuQGPDSOzjr1SNZasL2Ytu5cLhjjhNvRT6rTZoUdghQAZJ89NH3EZ
cfOhQG5t2/bOvp+TDe0Q3mfOK6O+1/IkSbhk+SeoMobNXXhy/njJ6fUoUcFmuZkKXyNpBxJ5dbD0
2C5UzbYnqTWUbAkTxgQ0BjLUH3JHDSaIeDWWUNV2Laxuj6YPDFLNPDu/EiTqLTb+0WBmz5oA5O/P
phcqUw/FDZXeE10RrVyYhnRfMD+T0JWNHBYYN0CnWHmZbxK9Eb4JlUC4SotBtYTdgnOxMzAQ9VUe
dDs21bU+Wcj/s5EASO0ScQSKdHqqX2+aUlnwPRgbcN7Sal2mQRIIax/gkPvzqqXHOn6VUXYZGosn
Q8Q+EK6rlTeONdJxCe5nbDvPOUargnAdH20BXNyeX3yY7Zqtht7gz/Yhd0NxFwT2pMqhD27XCbbu
V50/LLyU4YYaKKDAJP/Rn3G9Hmhqr5Ge1VmWYe0oLj71GkL404LHjbvIOvN+hboHPL5d3cFijgK2
H23sIL6YHx8AT3WkCryqm/sUYTJpYH/GZCz4C+XwS1A9UvQ+VNadm7eYLU3PPJqD4+JVXHFfIBna
GX8QqVRh9o1TzF1+B0GLvWjcF7kZHRBELOgqkoZbBWKa9dMZuVHQIoeCo3BaZcbvMZasXCacPk1c
Qh7Ic6SZe3eQQPNXpwLURtpWF5A0DLaZRiMLEtP/eFiB4DT2y1uKDl3Kc7YxCvJ/zu6YNXMDrv75
ZZG8kBjNeiME5yP9crePvFxMHiZzuNfaCShxMrxJXdTBNjv01VtEnaqHimUDLPEJFjBCoikKQZhu
j2TAz27WMcQYD35YEE7zxE3TMfXzk/1fvnQ9men0dU8upi/0451p/Pz8Yp+1z0tzF64lnNJEUkXv
8mY3/TiYqPYuqSHRYI4+JGs2mvBleonr5jCDuztLOgPtGGE4b+CLYcGFMKP+7VaPXggLEnFEOxdo
o2H4ySsJacmQiTl6sAeCZeZBd80HKD7HSr8mjJHly6kTIepXSL71x7a1Pz8JOCYSxnNxL09XD/L8
0iyLAoKtbv36Hui2oftuCqIDIJKmSJPr40VL/WNIByjwQPUKMqZ52ASTtsXUSYz3OsbImMFC5+nc
LzjxV6dosABOH2k8o3bMskkF+l7t95sxhiYHbT4ac4BrRnoWFApo5spv56as4hLt86ocwBSRRoMz
ozW7eS68nF+VsRDAsVDRvfVYrlakw+J8K9ERAUDqXqgZnXc6b9+lRodCEuiPdF13C6YfMSKsSYFw
aQ3KMawxcZpjlO9rGkU7GoP//6h0fPzGfclNdR+pNXcpRctDpNcGNq44dmHIjeI2I+uHFXxfxcWX
jInkPQ9Gz16nMHzOGDCHr+1wF7RJejD6NQYP2pOy4MrVKfk7l29ErpApZyF/zGKYC1Ra8n+l8fV5
GBfRIeLxH/iEThltdOWUmh2h40fBaU5pU7ZtIMt77vJzOrThBIbWz8c0XWE76/bx2HbwRrKIcSVf
RRIwl4/F0xv219Hjqhq54urd5aoUe0npce4+hFbxQKkJ6qCyZW7I/W87NttGM5/br+2AnEhjmAF0
jlBjUATBRr6Jo35sseEKUbnJDzu9mGX+ZGzVI/wi7VK8HPXvjZ7+upaJtn02iAqa6zu1OdYYDmmh
Reuv9Bmit9+sf0i3XfCz1B5lZ90bzqdkDcAqp5YXRfzlslC45dYEg/FL4fujXxBUOy82PAW7IIas
kkSnQbAHnZnI3U60DeN0/PxvDfE9+m8E0tNiH4E9nekT1Xg392OKr8HTe5lS2J4KE/Eb+rHLGwNA
9sMJ2I+tRZlhEjEBkMFYHjRj6UDfaduTa/CrWdOXKdoaWq+ehIYRkTvahPxZNkoey3Puk7nwsLiQ
MjP/Ohm40XF3Gt/VHP53HBzxSB3TDAPzOdBh8KiTjsG2/hqajjyWS+ciDD3JdpFLtfUGP5caG8/o
YjP7quPNccUa4Jh4orv7EWYyKHhH8F2vm5BTQsZgyoWSwf/MbC76rlkV6gXs/aDeL5v4B620ZnGj
TyFuVKfNmZQqr5m7Ad1vm/L8jeKHRM1VvL3dy/XsBIFhuPeMYioSOrGopS8G8c/fg78lhdfg7TBQ
+fe+OpwHsU7dMJErSR6OESBaFu1AOGPW2BZewI7zFZdC9jD9ceMYUtp3btj2xurNMw80u68OfKMs
JvsquttfQRlhk1bN+6c6kT3G80tNcJZ960Q8yvDnD54sXlgaTE7XRIrLo8uJY1ifpGHNbckuItiS
5GF1J7Ivaf37HfArBbFBvwHpNc34LJf/WEagF5Zqdi5Dk3HEXsNXQyOCdBhpfvokM6KtwiOj+gjz
/NeYb2JqYYvolZBfghZ/ICchEFpE2LS41Tpefi1zAQsCJkZh9ow1m3QCvyAzFDh5u5Yli1RrHf0H
+m3MwL5TJGC/ygYSoziIAFrQivlIGf0oZ3H7qqVlTSDve/GWBruT0T+dOmUUilrbKv3vPQBKCRqR
Ni51QkA9jLunZYgEbqdCIbAN5IijyQmb/e+8FXdFC2YEjJdntfBWEK9HWSdtqD36gudNKqVpH9bX
FCPwEQJX8plwpt6oNVr2BalHduFBvaoq5IhGT5v6xqj0whrHWVEMlIEpWzY5Prmd6pqhqvZ1CEKV
gdJvtaO35GqsLaKNh4h0GZBed3+9TtVdxNHXC766dHht5Bd0r4OHWRzIPtcOX4nmxicJdzsCeMrk
PUG+wa6AXaDr0xImjkPLc408f2NdIVpjj3XhhzuEV1yXXeWMWQ58jCd04kQrQ6cNqS28bILDoq5m
YMYZkY3y/0Xkp8T5BTV/zZtTUmvWnWL9w471pzP8oCa+fxFv8gQKip0FHobWpiSP73BRPvOn2HUB
OC+Z46/2rA5BDcMzQ7JNVEhQVcFYBheTU5iZ9uVoN1CNZ0D8P01Nh5akzUrgglKnUS7irEiHZoFs
c4L4oGMA09UKZhYdcsIVHr0JoE3Sk9qnWrfpUZXyQ0egh5533M1bCcL1mdOxSYGbHGLDFbYJWhIk
Aivyk2P2+oaCddppy1PB3y9ccX1/JX5rScgQXBeTlGvxW280MzqkxckWy5mh/i6raolR7rTYxgdM
SyzcAVYTt8M04nJjuTm74iZbEXtrlKrC/2dm/SHajCWrXqx+y3Gja0desbOAQOP3idVnMswaLify
tYVVymoJyj6INqqALO1uqEZ9FFTIT+fgxTNNuAJY0h1Kh42mKKP7pH6Odiped2Pp+LpnVc63HUHq
bX70aPpk7zk+jk81Kg+Rgxj/oOPn7/ew0EO/EPPtaUXc42yi92i8+dFqgzj+pnql1LLP/wtdxDy4
yoDCrwK4vBFKcR3ygxrKgzaIzxxf5diZhjyvFaZ9LBIcMoy9zLjWpoKbBvlnoAsihf+F7PVUmJYM
KmqUPWnL3zlY2Zhm5qGOlK+Ul0pqd5ybU/4sGPBiskkrUeEdIugjEpRfohJnRQgQEeB2XofUAScF
b81Gpi5ZeyVDrMcglMNr7dz6bdDbtS/quUYLBm0Z5C3iR+e04AAB3fkmaqbAO0u0hIoPA02iGGsZ
ChmUICyWh73qjdUJCGc5E+3bBHiXsAnaJfbsCfw4UBLqSQEcp82MCjq4mWwiF83AoKkSOR/n1QC5
9IOAFcrmdnpZ38bt0K5aLS1bRrnlgMnA/RXDBs2ZAj9n7+heGqOblyCmZzZQ
`protect end_protected
