��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z�����Y3�4&��-���"?����~[�Za�p����@t�<�l��i����V�"r���+9��}�E�-i�c��}V$��-��5�:<~�`�p���Y��ݍ�����3�B%N�b�#���d��;������������2���zff�*�������(�)q���"�`!,�Q���c�м!�k�I�x��5[���Vo��	�u�q̅<���>ZX;_��������r��RN�_!X��u:�Bj&j��ڱ��k(^��|�Nzwh���U��5$�������J����O�;o(�B����E��)��W�o�'�"<M��'�����9isb�渰D�|V֧�0w��	��Q��&�i�f���[����?��a�`�\H��a_*:��W��bY���g�$�hz@�� u�r�ޚh�{�g�cP-e&�x�N	60��M�+��m���i�p_�|���z�Q�\f-s^����w���`wR�m�I��{�vV�O�Q҇�F�Z�6�Z$8	����<�ϽK���T �W4�'��z�T�d���l�wWm[�nC:���q����V7�D=S�m+
��eXK��4��]�Z�����_�~��h&�\ac����z<E�����B[����=w����F����
H�2<��Ϳ6:�����#��0+�ucc?c5������8�Ped��!�g~y'֖�Zk�P����A�H�ZE�@y�i����a�M,|:�[V��a�~=I��6��*ē�@)�W�����uT����?�y�w��N�a �a�)2��������+JeE�P���D���K�v�qb�)I��A��q��j�症S=}���{>���c�t�������c�):��$��ԑ����RlWT�E��m��i}s�{#T�ϋ��&���.�Iҟ{�3��@p��<5s ���Mp���,h.ƲtUX�;�d���M������{�`,��dƝX�j=����p�"��g³�K�az�m
��u�G���A-����V��	�׿S43���9	ӐE@s�)�j��KG1�D�b:W�m���Xl�d)5�CX��������'�_��QR�;;u��_Kh*~��%�sEZ��=t�HH �oWbl�Wk�לdN�m�xԤ�	I���P?C(��F�mo���A_ض(��&Ӊf����)�i���Az91v�J&����b�Q�$y��#�4:bB�.��f�%Y�o$θ�n����3)9붻h6F�RڳC^� ^���9��[e�Jaz��?�n�ɚ	��J���J�u	���J���I��z�f�_��J'~�����OV�)|U��������C�3��{�ۖ��(����[&p�IDk�sn��7���%�������{�SѼ�T"Q-i�\ӫ\ք�xl��)p�H��@/YhM��N�f�(w��8�x��b�[�$nV��>
47 ݯ����W�D���漑���ߢnH2xl/�3��}j�ܯ&���B�����0�\?4�Pÿ�BE�^Ҵӛ������Rtӽ�(M�Yo��[{��Y԰,B�- �-�!c��@[��x���j�\��V~�U������9Wc�s� H��f�����	��w�����P_�2� G�����EA��W ���Ž3;+W;
>\Uz���aU���g�%�%s���2�.������H���֑�~]�G��kBTqr$�H�:j�����	��P'��:�,��� ,�9� �yg��C�t5�X�N����7<X%�[XvtWc�5����l���c&��i��ʤ�2���ݯ����������p��n���b�d,4o=��^�����7v(�!�=�4�֓0���0�Ӡ����B�����q�1�1Dj�0F� 4���`,#*,W,��@�r��sb"��c���gUe�2mϭ�րT?�o[:
�
%��>���n�ێW��+��m�25Jৠ�k�By1A����ܡ�L�� �7i�NuU���8� ���&���hT� ��9���1m�_y~d�|��a��b�׽<g�_G.'���/�A��h}�\d��KL��2�Ԧ�Ƨ�Ƿ��:ߨ���$Hn\�B��\��#��_L� ��=�amJ�H���T�v+.'u�b�ɬ��H)BD4�3����I �4�w�����>J6Na�&ӧz>�~,d_qu�%v���S�A��$jt�E@6��p��D���#2L KWj[�)�7�6ng�Y����L�y��!����e/�no�Yl��J(Xb��*����o�㜣r�D鍪���h��Vt��[0<m�D�ֶ�_g�R��̵L�
�gtY	@p/�����%#<�������W���Y�9tUg���7$u�a�u��d���UVk�@\&�����b�3l@���[�A��H����DQĐꄹb������'e;��k�A�5h�u��7�@��^�臲�KL��雮D��
ھ�V��E���Hc�:$i�"�<����p8�hg�h}��8}��|�k0)]����/����$8���ֺb?'��'hm�0L�b�Spo�J=m�"�U^�fj��#	�'�6��r��������W�+W��Ps(|=���O�|�C��u������P2����=Lu,�aύ�2n��)�՛��?�S,=Xm!9���-�7@VFQ9_D�EV�Q�[��L�����E�*}1�5�V�4n
�Ob�DJ�r�p�: {��VŔ�:UQB��&��/����:�c��0�Ibdz�+O�k#6�
��Mm�"7w<}�\�G+�2B����1�����|x�ͩ#s���w��cx��A���1A�qU��F���
C&��  ���$���0k�_Aq�N\��/;G`�5Cmۖ��	�!K�ФQ���,>����\��j7�_��i��{�a!3�ln�Z�/0� RE� 6́)��

B�O1�&��},e�=�� ���P��(�68R⼷��?��o��+�\�O&daצ�-л�l-�}i��r{�ʺ�tZZ�\d61��dh�ktR��;:q��8�^����D�<�Ʒm3��P�~ڴ�̣-]��R&���1�MQ���;�f�Q��-z1Z�3ú���U��YM�m^���㼉��)���W$R�'���9�q�XS�Id�M���I�����h|fHy��Ea�yJ���,x��<s���^6�4�G/�O�4;]�M��ک�0u*�j ��X�^T��m�HZ���?u�1�$^�[ՅB���t �g���T?��q�Z��E�"��AAХ�iLw.�	#��6jt&�X9�xU�����T�M�%��7������Q�\�&�"�)}���/y%
�X�}��#����3��^숨$��%ס0�!���^/�a��w*���p\���NH@͜o���'�԰@w~��˚� R�%�B����N�֜��`c}���%Q��2��� ���4��f�Al�slP�W��u>׭�2�kr�q�=�}#���_�P]�S��zc�Ns�M��\���u��\�vF�!F�Q uB��A������z����#�#}���$����A�Z���}��6��Pr��wf�;��Е���7\ %1� � �������%��<�_�����y�eS(2�te4u��|����{�;p ����Q7�U���|�E5���T&�Z�_�"�S�nAj^�H[8��we� �\�#f��t6r0pmO5�>�j�m}a�+v�E�?T���q�R&�����E��k�|�4���T�
	h��~����
�2fA����������Ƹ�.Ɵ�<M��T �Tۓ �_S3@f������`�s�`_�5�)��cC����b�CV��0���3��R+Ak�xW2�K���\k*+��a5Vؽ��<�����;K�Ş�W��Ϩ�G����y���l$�ψ�Ky��'�ڴ{;K���<�	GUUz�na"�Ć�z��@gOnB��-ܞΐq ��}�:e=%�Xb>�#�]�|�d���f���'�M&��WI\n�_q�W�G���Ery�$^�9뭷e�X��
~��m�/�v�Y�/ey^�=ze��~rRxI��e�K6�Z�K��BG^RY��Zd���ۜDBz���'<t�6ؙ8�0kV��}� ��g�MG�&C*hu�����$.� .@�9��`w;�}�뱐��`I;4F'D��)-�4�,v�([A�i������d�p�z�u�E�_"�^�\�#�(�6"�+ʯ�w��a����ѷD���"o�[��(��S�#J�L�4���xWhА�t�N���3"��d�t�~��P�w��K�72�D�/(���X��gN눻deUF�}���&�}�������s�+ȶ�����g�[ҺtEWL|�]�����Ɔ��#�1`�n$v؇�#�՗¾�.�K!T���'�-$���|.u'�m� �GzL?���雞tatg3�Exw�&%Q���%�?�3�}�}q�'Ɠ����C�(ڳ��J)��X��?{F�x:L������7[N�s`�d�mnc���v��������9�{��3! �`�.3��c]�,�n����C�%9�9܆�ށW4�E��úq�)��T�k/�*u�F�ᝍ˜b
8���Ij
�Gx37��bTC�p���g���D�g:�4�7�������ǒ��dm�r_�ĢӒ�aV�~�n��~�Ǐ�T�4�':�����v_0�:���l����J�S�RωD��L��Zk�AB�=��Ţ2�%�M��X��.x�JO�ཛྷ}ӛ��������!L5�U���o����ҕ����p'}{�5��	h���I�J���*9�E�4p���O�ܜ�BҨ�ef7S#�C��8k��@��A��ϟ�?\�����w ���\<)�OJ[�ˑ�����RS*�s]�� �&iPу+$+9�3~�)��)*|E�[z�.���W�g~����^n�x����I0��?�.rk�D��#.�(n��һ�yf��*��O�X���9a��C@_�1Ж#Za�4�^���IR�T�������i�EmZ+��Tڈ�u��n�V��Iq�!�giBhB VX-�6���Ng�x�����	��D�}M�SgZ�<3������$
�r�����\���
\�D�����;�gX�0C�ѭd�f�:m�<(�s�� �)%�ԡ�  �����=�=��_B��5צ.Ah�-�}���� AK�x��+�A`�mG�V��"���s-��
��#_����n�� ܐ�4�
�ajs�:D���r�]�9N�:x?9�,P�wʑ�!z��gm�����/��~���!�=����?�/?q�
^�"h~FV��%F}^�P\��k~��D]�ff���T�倸I���g_�}��|��9�lS�IƦ�"��~q
{A��h�#`�����,��42[�=��e�A9��UD(��ёI������E��X�c�Eޜ����Q��@��6e�=�������K|�3Tq�2�.���3��%E{�+�
߁7��`��������N��D4����󤀁�
kp������5���
Cy��м��|��L�<�С��]�7A��
��uÁ��` ��_�D�xL���O�5�+uy�Pm �]	���i�*�*�����:�w��%e+�'i�(��a���@<�����m�P�/�Q��<�k�?tɺ��I�s��4��^��H�xug���9�-f��?��੾�z�X�Tc�_B���c�����}�w�CՍV�ZU��ѣf~�%��<1�͐B+<�y)$��t'"�Y���8�L8�N�����ŤJ�|��{���R��>|(bI�Uvm)ޗsG)�j�a�[ �Mo��υ/e/!�?�G���cU���xa�T�_��Y߉#�:��WyA��<�x�4YVR��P?4BE}�q�"�L�W���
��'�c�y��!Y���\�֯��<�v��&�)�\��}�.�t�/A��9��04�Ɏ�z���dJ�0'�����@�n�����I�߮�[��L�{j��7,p�_��9������YG���6�0GI��Bg�U�0�_GA��nòԫbh�7o'y�Թ
e�=�Z}��ӄ7���9��`�@҅�F���DK� �s��Y-���S!���~3/��*�
9��E즍��[E�~�4�:V����nK=�y�,3[ĩ�bL���^9�@���(����0.�伨<��~���1�k���������0`(��%�b
�����{	�����ɫ�a�f������ܲ���F>%�{��o�F#@�:��ن��.�-B 3u�癤�8<d%8jG��ꏀ��L���`�{��s4>0����YՋ�<��ؐM�iܽ�|����Q�<�C��_�BZbbOG�� �he:���H }	�?ѱ��M�5�����p2Ix2�Gi�m!Q-�Y�첢KF+��9��r���G��%�l��z�fl_dU/d2z�j����S`��11/��Lq�mw�0	�4�H��d"Ft�?�����d>U�zQ��v�o���I�Ֆ�R?�IĿ��4��^��Fq�8V�P�%,����礞�� �����~���kp
��9�ӫl�W1䏹���K�A��z���N����"S�u�;��/"�+b5��?���kqX/�=R߾����|Zf�ETg������*x��	��L5<�LC�Y�m��bu�����!���Z���q�1��l�-�����-����YQ����*8�D�!�\z2���Z��H 1�Xo�C�^`�"����ӺIT�b�f����
�iۇ��-%�B��d��[���X+ycEsό�K��*ڥЩt��1��|��#.&�|�'L���_{;&9r�I9�u�fEcf�ֹ�}2 �q  >�m7}\áu��^^�q�*3D��o��8�O�+��h�����
]N�|�n���cTQ�$7�+wT�������
�r8dޚ�"�[�>����,�F�By�rۭ��j��o���ދ;�\^�]����=����s�?�����֙���HpB.��_!�sG�.�c�5�_g�`�fF�r8e��C5��^:2�^~�#_�O��ғ+tI�etI,����e�V�_�f����#N��α��#��"��/��%D@`���������__Q�Ǳ����Oek�i��X�~c��irI3Pw�(Zqj��"gz��򧎲��K�ME��H��BJ��)�bo����Cfv�^H�-`��ʩ�=�]�2�*� �wRy�T>�C���_�uJT80J���0F��WHE,��{R+����_�/:��`"�ɂ���5��j誢��~=ڛk����͐�:LQ�9�%��͑�N3P�(w���L�)���b|�wY�Ս�|��V�;��7�V䍵+��{٥�ٌ@_�堑Z/�U��u�U� �,b>lv
$+�4��!d�lR�˹���$.�wH���m�N��s)���/�H��"�~�eC/1w�\W��L!ԱwZ(a�ݸ	��37i�����+��n	KS�8C��2(�l��L����J�ȝ�1a�~MX�Ε������Bv���b�NC��m�#�gJ0~��s�C�[VQ����`p�ބ[n6Hi3����wαD�H x����m�P�z6����5�u�cr�(=�$�ZWb�&�;�h��U�2!֓���{�pΕ/&�|s�D���ެV�H�H��N�&����,a�+�FM1�;��(8w&+��^{�;���~��<�^+nS,���ÝU�XdQЖm�I�#ຫ��F�C��8�q,��%f/^��fJl7-��'����[Zh�:hd����5c*����cp:�
�����8�7W��ǳ�f��q?@Y�{o��7��2ۊ��P��wn���9@Ҩo�*˹˙1f�O��Ld�bS��60�vV\6��\�^�[P������@>y�
�c�З����a�Y b�AY,h���T��A&L�?������ͱ�J]�~��^Aݜ��}����k�N�q��iE����\��>q&ǌ/�����3�4���j٫)q������?��L���ڜc�GZ$V��]eC���_����.8�V ��N�����4_�6Lu!�Ȯ�s�5ͩ��ӂ������/Y�Y;����r��wrf5x9r�"��gS.���M?�a�V���!O����1���S��o��?�|4��q[���n� Ym��^Sq���R��j-oj= �SΘ�)<BH�����ɳӿ�ڗ+�:�RE�bRYH%�oP�4xT����?<_m��k��;H�P� %5�i��l�m��%���w��:*u�$S߸��[a�]���o5F�˔7m�r������y����I��ስ�&#Ц�zWV��UL����C7�;�juV7�+����g~w�P�kX��O��X�ݬՀLv���\��$�P���t�R��b�ϳS�(lܹ�b�o�D]�~+a�f0r"'Vl���.9�_��Ur��C ��6�G��GV�l�Z��F�i|ѵ�-��'&de]Ƒ7-�3�)�^��߀jOU���4�>�n��ϓ�K���a�"���G�i�,\3�:����ȤߝaӵV�d;��,X	���Hxo����am��b��S?o��F]іKk�����۶�&:�JS� eGāa�d�� �I��J�Lp	&��"r�-e�,pb�mAF����tV.�I��l�:Qi6͟�>�~����I���s.2W�W3���$��[-��vĲ9l��D��E�j�7�QR���?���f����a���Z�G�Y�'*SNGH9:�$�c�N�َt����3G�kE ���hͺ,(U9ڹ�6��B��a����:��m�{�z~�S|��l4*&B�"A�w��HNd� �:�Q85���E&�{"��%}h�;��#?�����
��f�-�DrG�	� Z���ߣ^��Sa_��fE[�����&��̪-�����Y��n�b��ן ���8X%Y���E!}���)�lg��Y��x��b���u�F_�(���^��m����]���Q�b� �w=7U�&��{b&�Z�S�E��/��`�Y��AMUs/_��q��v�G�{�Eȍ��ω� _�s���,E���ݹQ����gK�WOa���tc����&h,	G�y_��șr�Wj�����u��ΝXS�4<1�h�L3O'|c����E_�8EY�Z��nS��,9���
u:�Wr
�f�b�4�w�x�!�	��"}ׇ�_j��jF��״6��B:ZKU�aZ�i2b���x�#fn�q���*�e�(Ab1�%�5�~d��ظ�!�Ve�㸦xK��w���4)AY���N�#Lh;�"
���`��s�?��4ˤ��E�U����e��0u,�q�ڲ���ܨn��U�^�ݔ����}]kܩ6�:�Z��2;O2�y�k�Q-q���w�q�Ϣg�%��X�b�>�,�'~ĳ-����B����mLM��������Ҳ��=Q��-��@�����0}���ﲝ8���A%+��{�%���l��_����N�'��|XP�]���Вpk'�O�6�����Z<���[���܂8L��E<6lOE�����H��C/��m�v-����l{wԭl�%���WВ�55��Ԃ�oZ~=� ��O@B�ğK!�p��4/��ޏĄR�,A���k�&�!���2�\rq��	§Hغ��@�b~dEZ�19��VUo hS���.?\���ű�U�n#�m%��ӌ��,���ok.���L��嵿��t�G�)����F��Iq�W��^-1�aI���"z0so�b�;r����񐅒$|
��EU�R�O��.����I�� P��4���~��a�Ы�ռ���6BA(�ua���	2^��
����=62��Lz��`����a>9�hw����Pi�G�-�}��X��!B	7�Y@1L�d�[|��P�i��$Ll}L���Y>�C��2(����H��lc�ޮ�/�10���e��ܭ�{j�q�nB�i��Id
h�r=��?ʘMP�:���y�S+���v�&��@�
"(vV6�4Ƹ�x�d�{H�ᶵV��M	`x2~Z����S�*}6�B�zg�&ǵ�8�4�h]�
�5���E"�B��ʆ߲�<w�"�C\'�{�gR�b��t�E��w�d��]F�p�n_l����Ch
t0�J���iw]Bl0�(��_��Rq< �Bznu�H���D�����?�� ���vJ�B�w%g�1V��Tu�a:!��Ȇ%�7Ho�+����s=C�Lay�镬M_q��eh�e����V�w���ʬsu�;�b�E D�K�����j�j���W�d~����h��"�~NO�%�j8��`|?�`��
���֕}����2gM��6�ge�d���b�������ax�a)E94\���,��a�{��1����I_~��-�_��.��C_�@�p�,��~^�j
�7��ލl�/�8�6�Ԋcu�;���4��C�H�v�D����t�pn�[H{�i��ʐ�!�3��R�(��\�Y��Հ��F���:Ǘ�]A.x�F&\�>�`1|��4R��s�(��{��N�T�W�
���s����I���S�M����L�(�(��ں�d�ŻO��H�&=�y;�	h�"�Jذblb"�]�Y��
���c��muR���r�
u�5���T�;Q�!⦄�����a�`t�2��m"����p~{[;`�����Ġb"��4�������a������e��B�i�{����?�v$A��~W!�2s�ϭ�[��l�^S����j�ʷ�C��"#GM̟�06gҴ�^f�E��
�@e�sj#ę��P�G�$�)I�_�*An;~X�n/�W9�ɉ�T�c���V�nQ���~�+��R��{�v�pU�C�8�/�,�R�T�8�������6�Hf�V)�~�0�즉Eiֺ0��8�#.\�����W���*���{�f�ӹ����z4^`�焟�T�y�?��<�� �ΐW�sG�㚯r��:eP�/ۭY��\���4��q�Ӗ���2� � "�?��y���6�+$VC�wZfBJ$�L�Y"�P��� acOk�4�3����z\N�|R_l) �@v�5W�@7�����O�_�����$��i��
����$��`��/bD��x����D(����#*��6As0���~���k���D�c�pt��ߞ�A�g/����1���nf	.�l!AU�YՀ��2��M�#zgS�� ��g��Ή�Na�q 7ߘ�n�D_�֡�;���ւ'��Mj������	܀[i��`)����o.Մ3�iQ`h�2���rSK'��CtKq�@���~���FCj�M*�NQ1���ax>^�_��Or`�
� uvXz܏(��{-���n�(W��޸G�|T<z���/m��@hCZ��iI�׃�C���q��:�Մ���6���3��8�,����ŗ"�x^[p���l,n�����xޯ�"L���fm�k�`��ap����ΙZؔ4���X��MI^�5���c�S�ˀR�����DBu�Ӭ�����"���Tt�AH������\B��~9����g�=po��Ϸ��N�y(�;A<B}D`s�A�����lP��G�"[��O0�ƖH|�nX��`������ں8�(B�l��I+\�q���f�� ������A�n����(D�E(��.��h��/����'�3�t$h���c_X��������E�;i���v~K�AP�f˃XdH�(����E���*���n�R��E���:L�-��"�̼�X^<ӱ���G���2��tX�#�e:����93ASMu��枰\�����-j�7��w�	inȖ$�T��C�|c,�xD�� 2(^�ڬ"$�j'<�\�V��QS�wzX��@���H�Z�rE&��ک�Hjﾁ�b�H�I<�3��=��Q�+/�O���F�l�guFQ�&J���Z]:�κ�?�]-PU�E����7���»��K�p뉅UZ2���<j��0N�tG��V@����(0M�I�er|�u�t��u�Ӻ��=��1^�N��ӗ��Z|[��mIm�9Wf�+c����b��[Zǭ�c�/��෉�a�	Ly>B~"�q�n����q]錅���f�������>�h��rށ���%8N�LE�w��"`��w#��E�7v�@C�'M;E�N��T]l���Ck�e��;rƐJ
u�Y(8�`�3�<]S����>����|nǐj��O�N32�$R	��sx03�g=��lv�m���Vq�]���������\�(������?!{vr_��-��BC4��R���`�m��Jl��%#�- V����Mz@9e]}q��6ަ߻�6z74��,.�Ka|b>�ޠ<�w����	;k.����x`��k5����ëa�/ �g
�dh���n���oį�rHV ,�l�y�d݊�))��*󗂖���3���Ϯ��`\�ן����]wxj78o�1W�O��q�P�C�Hra/7�k��.�p=�N�\�U+o�����(cbYr�e�e�9��<��
1o�!8�y�N_`�qQ[Y�J��ډMΒb`ES-]����z
��:�|���U�v�Gzak��i�:�Q��=p�झv#c:�!�O��zO7�������:�qK�� �V���;�T��0�8r��u�d����@[���դn=�)�	�e��4@����:���߉�B- ْ���/��L`<4S�}IB�X��Q֌�>}\���<A?��X(Зd9���	�:����o�oxTw%p@Yn��rx幘�M`k{\�>��S�:*�{(��7�¹Uq��uaC0� kE�����fm�=�>� �&�QA
���k'k(UR�a�s���[E2"���af�q|�ƪ:$�P8��KA��ù�,�&E�x�M2��ˑAT$��Þ2<��b� p���O<lH'��h���ȭ�FɃEP  ���Q�t�Q�m�́MUh�%�Kͧ|��ڄ����gb(2����E�	���S�=��-��4����y�����k���!��~�l�v?�%���\��N��p�Pǂ�i\���>���G;	���
�,r���1�|��
��|ʹ��2 �kd�Wz˃��~A[��ֿ��Li�Hm�x1 h<�o��'��C8�b2��٥%�G�>�T�b�Ϭֵ)Ћ��W�D�u���p#`գ�Y]2�̨�[O��e���M�ZNni*Ի��n����}�m�+�?\8�B쁭�jE�~@���M����J��L�I-F�œGA2T��,���YZ'R~̛j�C��3��8�=�H�y t
]q#%9��я��!�R�E�K"�(�p�*�(/��0�oD��སSw\8�	��#��](=��.�Wت}1����+�BL7��՝Tc��|ѣV���
���}�K���4��fW���P
W��)0��L>u��0�#�h8M^s��;�M�i��5KҤ�|�>����krn�=���4��&"��=��I����Sf�"O��� .4W����S��CD�M�G�)y��V��S��Ր��E�Kom�0�Xu���tΎ���YR��j�	��h�!%�nm��P��c��a��Y��L���o�F��B��~Dܷ:��>k|��4��=�K�#)NeL���ԃ��f�����<������$g���[�4�����؁���iҦF�����)|��p��tܔz
;�0c��^�5�l�}��2��� J��N�mع�n���C�ǜv�@9]1�eD����sY��+��NA`!p��GQ�5�[�s��$-��cQ��(����a֘��D�E�c��L��|�J�.���ۜ��r�q����(+�E1̜T�|b<ή��q�%�*����12|��p0���:O#o��R���Q�ǜ?���7kr��{ʏy/�K�]����]m�Յ$۱ʖ�RY��٥���t=����!ՠJ�c���#�X��[�}��NC��J�3���h�^q~����N�K,�T���
���[J�c�직�;�閩(/���Vq�m���� a
����z�6@m����RHH���0�%�NP��薹c��Cō��pH�y)�Y�@��h���q(q�� "E��Bgw#��/�!;����XnW8#��rk7Ԡ+�<Ղ�2�fWs���cΡ�{��o:p8�Ԛu�2Ch0�����n[4L�L��+>�2�qК����4��gW�Z\��/�-�qi��.��EC]�q��"��cc�,Oh���ӯ���u�����+�H�ݚL���.O�X+�'s[�g&t:�#
[�GVg�.�kP�������/K���~�#B���t���k�9�$�����	���_(h��rOU띷z�cS����.!�5�4�3����c����)W�񁷠�$�Gz�����n�{�˖,U���9�Ʉ���V;�s�@CC;���w��L�͡�̪��U��ώ���DsNsW�ɩ��c��~ȝ"��pFA�:/C����P�+L� `�'7/�,�V�uMB]U��������8;�A�֗J-]�}w��<~�;����H��^Y�o=��No���gv
��޸+�ِE�sj1:��6>b��a����ϳ��e��@YAk(����Nh�����]ݐs߂��,7��ٺ~��C�+��z�6�<��ұ��SG�]D�0,��w�8�-��I�d��8Pa����\��(
X��l�I���yޭCwPIo�C�=�zZZ����������q�K���Fiz����݉����}TxWi7C��5(����f9�Q֜H0s�os�%��}���ʉѨ�28�M���M�d��ܤ�ۃw8-�켜��!v"��%��_>���l�MJW��>�i�f��嚑t��P�"� ���҉�g~%m��'���\���-i�{��g�QN>�ߴQ�Jw=��`�����!�f��I~���[���d_I��z��-ҝ��R��YO��49	vLS3i�y2�!�4��@c=�[0i�6��S�;\*	�v�R��R4^�u���U�.���m��jL*�nJ���R���G�<��u�-�l��R�ZȤ��W)�q���©|Bg5x�$��Dfی� �X��Zc���C8Y3V�}�K��'h5���F�Ƶ"YX����6�-%��kb�Ї���ὀ6H����-�-�2Uf���-*p���߽pՔxZ*[�=���DS�dζQ8(:&��4T��+5��1P�K�z��ԺA4�4��#���Pa�Ҵ�~\WA�K?n��>�A3��:�8�!��b�#[y��q��C�ܗ9=�c����;�Uެ�����n