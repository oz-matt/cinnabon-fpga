-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
YYmdmjpbguTChMtF1zS+kqCBIpihg7Pgh68WkDdPuaS39uc6ZE2n+kchMAYwXC3DYRiPJPtQp766
rywwBIL6oU5zSgEwprmC/dUF8n4PbBA23zH5E2Cuk0ImuM7lKgybezFlI4K2pnqi0Leod9jc/cmL
Ke5gCpkTaPlsm4R3hQsyyLtKkEHWcemt0RfpnpF1vN1CBL0xlYunfWq+lOjFAdvQSx1AEQuFRvMA
6y8YRu9Vi/edeUPpB1iSc8gyu9/MST27tCbxmIee7pA9KOSS9XHeyIeFtf12gJgUdP1Nvgtazo67
aCepxigx5BLjAasPrFhXbt/ITqnKwMB6xI3MFQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 12384)
`protect data_block
AxtEZcbbsNCJJ27HlO338ExEYy/1+8HKdUSO0Y4KfxXmiTxYVdCl+xmqEz+U5xMo25nTwOhSmWi5
q2suKHQ1/2hF/EzedTSotMWCTHPzgmTRmchgqXTcoU3bGJ+0D+mPLPk9Yav24rFpu8qO3mqLXSby
l5dyC8KX1IgLhV5QNB2y/Ii6NnochFpT2h3zle/nQNRswYU86llOjzSTUSGF7zM/aOarwiJKQjhZ
+gLgn3HfDxUF2pF1HoooJcs/A3LMPrLJLwmiafutIWZqevMYJv8az7a3dIzifikUDI+lK7aupMNr
rLCJIop8TDWc0Ie2ANVy/vcxplL/lPEUtR4SzS4zSefb9MKhGcbC/uiXPvkZkgF7MXOJG+rYMnPb
YlXZIe6KlF5rOWaUSQn5Vs0nO9OlzT/xbkMEkaUl8sg77m7xyhMv8KyHmYDzSpHv5PKQLzVpm+YX
3HemfILoeY4MMKWdW8NONYyxGcPZ7iLQrIDY2U8bOopXByPw58kwl50IUbNM7hBnkUCO1ZXwojIB
mqNgdVbWpFtTFBn/mcQBjuTbVwBG2y75miQE1QM/auGZebM8rh8qwrJNGP+vnoWYT+c2Nq7mhsOB
8E3YOw4nYbskPISL0JlXjcfwufM7eMoHsyoLt44qOjqRgT0CMnvAlH65TDDAm1021jo06gCOFKxZ
yrTK2P4t3RnOEkB01So6nALPdDvdRNjt3OqdbONgpGlRSms7TSdW1Zv1/bDclmCJeXyGjbHIEieN
SIifgTK6l+nbpkQOuWHNg/R1uYU6p3Z6i+TqLZgM6s4wE4Ih336/K8DTvGZlJlaKk8DV+N+64DD3
f6I0xH4XKHeGJ3BXJA+5Eds4vGA8RLDnjnF3pY9FDl6bBdFmsMe5UNRyif7IyF0xLh0TksAxRO71
Xzd3r0Zu2oZbdvQvmGPJ//+DBf5HoksKYs6+YnTB46+Ltvo8xI7PgJN6/WTeUE6K2tQ3VNpFuRbF
llbDzsr6Bqz/rddZwYCWz/YLjfoe3LIs4Fj86IExQ8NYhKStvFGVaxMCrNS5zoPdKDIptMg2OnFV
xm1TrXNoySJgVoUHWNqsA6gl9kjue8fj+im8ELwJ+ba6fz246Cw5oM6ElnzHixksDYXw7mmZnu1W
z7tjudsM2900hjIe1dp5uPaKUeuTAjfAjPiN7Nc5EHBImeUgD6IZx8whfEs3fUVmi0GryJ4wVev8
7gGRxUM9mF3hIuiVUs1KDtOitTdMv6BpqWvxuLmEd5QiZ93neDd4PNpj8PT1Itn0N58KLEa3UgJM
CI8m8DnVQ07OFIF3aU88bKHfzd4aBCYnqII0YVMfqJSOl6DV1jt1E91Pv7YF5zqEVcmTlFCG1pQ0
0RYKoevkBETwEx3J0pvzWNRYrdVqgBQq6xR+1drcGXvn3jyKbh8Jyso6IUag3UzOJAj8VgQuA+E3
aIkUOYzf/KgafZ1HAyfdMUk68DvpfLVnFJK4UL8a412OCixXh68ZBF1IGENL4/QJEc+Mx3TU5PNZ
aulfjt2B62WtFyKMATV2dCAEmBTngtDgS+sb7QWgH9rYvoUFqoL6jLv6k4SIialJ+pl/x6CupKLb
C5MdAF1TDVmmgzQPc6L4MPYOmwsISXrS1+SDG/GUULoZP456KRiy0D2jyGuDuG/sU6YH29aCRcH5
QaAwTme7AEQHa7Ce/sTh21txSbUMt/v7tuTgRmRHTl9ccReNUXjo/eqxdpaQpkXSEypNj2rEsHYh
uTQ5bnQD8hgzvN27PTBCsOZHytTBmIVDyyd2892zlSjN2f1L3uPVjsknBqWlwinWmq3oxmokRb4i
FMvQMHKR+Xg6Cy+jhFfpjLrxTY/9WzXn+UjT2Y644liu+cXPoeZN2T0seS7J35tLTeV6ZqI0nSAG
ExR7lkX/PSsa42pE4BauSQTC2wXIPXcbszG1gfRx4IHvO40Y2mEEDAMKenHYzHE7apt0YcLPbsfp
kMWtSfHhqapI/I95M6BHXaPZ4a6STVwK24g3WxU+E9FlepziuxVtbxuK6NNqxHNfMivwQXM6lXCN
CmsyLrXA2u7zpHiHUGi4l4UZq/WKQ9yF+ZdbCuz15M/1C+U6zg0Y58g2jnCsZAQbeJdvgaoMO66H
aJliatdXLTtAw/9YVOHILHcr0nDPMq2HbeCVfFLNtZ19SknLJ1M0K/gvVupAtqayEM3N0KTTAR/K
dzBHw4e6wXiRX4NM3noV1FY301Mw2Dpj3Y7QTDPzeyrvDiTe9nw5wc7syJ7LSmXLO4bntygm0DyZ
VXFDfG7rpKNGIaNZ8SXwoAYLTqUUdB85RMyTtDZAP12jsksofjAysWngKwPX5Kb5bTSb6gsEPUlP
vlgIesBEi+4WDkjpQr1bP6lkRkXcgtz66G1Kmp4fOQBag/nuI1wrQ/9zo1jAY3sHcblypqF3LDjQ
TbgWiTuDUCBk2HAmMYahGE9Dmy/aZvrYwxA6Zwr6JttTtBa++4XGol0SPyV9jJcLyExt+zMS6KhQ
5NxQ+7MwrtywWSM+OP0rLwT+XRrPZR5NbzWP0vdf9V2xMhbuLFiPi0UCPMb8w3C6gGZLPHGQ+YpB
yTI3yd/HgbLtb3gx7tJ2eI+FOdtJ+fwpsQJDzN0VtyNvzQrzsXendpg2oZ2GDq8ud+ACsTZt1U++
Tfk+0127uZI4KOC4nzGvYegkzhjURkonSHtyyB32Uzap1miRoOCv4dJz5cE6zg+y1a2hxCnMi9Uf
YueV+v9lFcjfHyvtoOvJrzdGAQwdUnD/RZCb0I4y0nGQHoXGFKPizwwu6jY7zdViP9m07/Cm1sbj
bXjSJWku7oyH24hADSs2DNK5/Yj7+8yUO0Xa1Dgd/P00eh0ObrwMA+pOhKbqNA+vH8h3esrkLR9y
AvUb5uwysFjZMu1m4hVf2KM5e+cXyFfGvde9SPM9oACmP+GWPE2YXzWRTqjBg6brpP9O9rvzmIcF
rqZCU4Lkf+4gUTGfMvU43RoEl7BRKdhn3tw+bWUL22JSkinm8dAnSCRIBYx8ZeY5A+nfkn04BbNJ
Ni/q40JWXTzF2G6QXY4qL0He4Ozn1TwHqHIJaLE76V6W6TjQ76GMHFU8shhtU4xzyaD3T89AnnnC
JV8GCw1IHf4sCfplxktQHjsewC35D59dKRDxFHuptq8voF67oy0Gjh+ILm2vs9ccdXRlTfGUjRxV
CaYNLlYB+WHPlr6nCxN0SALIxiZVA+k6ybBvAliiwKmryZsTPSQkk28t8fOcH3vWAG+eCGVuosCx
JGm1ZB4JpGfuAYEHPdqKREM0fcNV5MsdCQ1yf8QVC3P4vE34aKcI2eTzK4oALBenSzlVVA1XVuVF
V4PjUNLjw+sfb6xhHWaxvRFzcvwEIerJ0m+5SGCyX3uTYup77gxFN9otUMcEGkFV8LKvx89Czt+y
/q4HXOvoSSIK1JjAYPzMwdxT3oarWIZDV2H+Sdtr3VacfCl4hyBqIfgd845cqDxx2gnuBb6Piwqt
iuMFHNlsk0FXlnlX9llddOlN30Hscart6orKhLazgOKrBkugg6iCPSdr9AsmunHlQJuAmObZdoNJ
c6/M1YWwPbxuSn015xjzU6k9lzn/azKrn31/8YIFxYk7WSuEEycN8VBru1O728UYysKGMWgjZF5H
1rlFCRgY9zFffuP+NUDPRj2GFrSrPvxAQ8veu7zahAk7vyz96TweZP4fssIt5rJb4BUZX+dny/7A
QT3DsSCsYHc/smqpqIMVOqOEFv48OjExBNIzMcUsdcGjjcMuJBPvXgctl7N86OfPi9cq99dPY+s+
WgsYkbsbtMXhq6c/6WwKZ2+C2CdHafiFRGTtiNtNCdS7d6+5Sy8xS9aXvgQJX82shoAx/+EIDyMD
d44NIDyG9TJAfXAzHbtgDDa1sRQTDEpz2gpnUuC2phDNQ5hrP0vPy9gwRaHSra5RFfZs1HTt1iMo
Ywf6mgqBosuQ4WFsuuKLqxJcTPBIgrlX5JKao9hX34dyetwW+uxTrCqOob4JYz03Msrf5BbJpewo
Lv6t4/STE7EcecN6j1MdfTMz1IdaGGfML8sEuXFkZZArDzRdw3wSQMbNkmhQurBsKaiO/dqVzeD6
cX9U3mzh6JjXl0jKWopkChLgIRCDW4LrjIOOmsu4PIuHvz6ry/BVloScByBMLRdi86IB3Fs8kN1o
32N5QorFY/vUCj3zgT3/5GvFZreCO0eXlpdJ/ufB6VRsnmXz42U7XHyMGWHjOrJnxkQmuwJx60cS
COD4N0uRbb6cZl869CFpOrcbJAoT7dsj5nxGRz/kYQBCS2dBdcqTHBKWLITeNudK59fcJAJMtIue
EgXKsZP08G+l/rQwj2lWM3n5AUCJIEtNDOjQbHgHwsAL6lS0W8KQE3yh1000BRlCv8BHar+JRIZq
AXCjMdWN9bwyO4iSiEZpj/jOsJzS/YPagIjzzytKJpULla9xROXtfOw2vI5uUnWhxw8EuVIcU0g7
CGtLuVWhOgxGNR/3tVS+Vgn38BNfj8TzU7NSxW7e5lEKfROi14VYRk8w2lcuKr2V511lGRaNv8mG
XZO7bhhBOkRFPgtwcSDwuNqAqwZJB/DPnlkZHpP7wJa+aTpog/xRz9bucWUz/vShQgQ8r8TXB364
NwBI2GpXY0PRorNtjOO+XKQAQDyIT5bFWBw2frbyBGZPdLqWRPO77Rq7gV4VgH1jKlwUe3AEGf02
6nS5QwThTPjmQW4NMvDHcL6S8+9LkzrEd8DisM+4G1goNjKigz+H8SFWg3BaTo2IX8NFjSvNjJpA
bkASqaLH2d/gBhytPk96nrJw1oeI44Ehqzdd1EGPGyzbdvQPvoNIPWViQmNx2R7Tkz1rl/wuKP4M
t5dcOVJ3N+l3De1wwdQ/R2s2dbw9S9pbHw3L7Ur+vCz6dZLHXo7/Vp9loeHPKNLuXXw14edojPm3
Bx8cSErOE1deamDDJlDKyB72kriKLsqFo5KfONAeJpQEyFb7IjWWjQsK4+4xkvqGCW5G42ioYrZo
S+Z3+/CylDlC/FwjBH1X1+hTN7g8FI2dYY2ky6LwlxgZ9wQ8IDjM4X5q8SU6gdhWMqwYjzZSzWxO
/+0TLQzH7Uot2vAC3uqnrOPklmT7Q48D0fVksnhWdWIN1tRMkGKlFAaBU8X54BEkqtrIud6TIHL6
l9ASSSHasadISVfwEMabDewc2zx/ISxgXBXFSD3uJxTqljlLyexdF3tM60fcUygO/befmT9G7gsG
2grQiNF389N+Pv3c/QAmy7bG3hf2esJo0TlcrCTBKHkWVL0QHTUHeDVo62k0Bf98BzsQsIaMO+EE
fivGKQ5RaGXMq+3xM4Y7xy4LG1z44PKg4siRaoSj1cK7s/cf3kPKgdSksc2keNZCise7ofoYf1gk
nh1H+JxGt3sY+oUNPY1V1sYrkrWxmu+9Kuk6A5PbDqAidy3y5zemItMsweJw+3KcHxzPRPmAEm8O
pT5nGVi9eFhlGqGAObi1009HLYe0q4Kc2t0Vcuw8VyEiGUDJXDFJZ2iOv84otaGYzQ3D4EzvlkAv
EXWnZJC4PxEXmNzjs5+BY7K0Z92jxO2d5B3Qz16BOfvvmEwrYVmPF1m44mKdFrzh0g5r0r8dkQuH
FmJd2i9X7QIhFqVxVyOl7scmiNWXavQNVP26keq63CSLqES4FWpm7xjN4uGRqCHjSnMAOKeZegPM
0ME7IacN8w6cX6/INuqft+Ry4f+h9vaVUB56N5NpWfemdKR7IR0nB22AHE0NF8Xe32En2Mc73Xix
V28E2bf3j4hlJ6gHh7k1akDfg/LrsecHgQmRWXxpRZtSLP+CMP+4S1ANBLQLiWnIXSrILMxf2RpZ
hKKtD3ePmar/M0m5ZgTQ7AwmiLa9/Krx/Ig1Gh+XvsC2tJJgdBO6iAowQj38PVfQmA6A8tq+jnLz
OnhE4evZ5gkVaWVxerZXe54iA9MQEiQtvOajLO81lkH2YVyuoO+odIUjZjAXNXcLhoCx0Otw9cZu
8R/n0ydvC9wdKX/JzPLtwD663cOxnkplF7WuJcPvkMhVqi1j8W2QCZUOJxEkJNHZ9pC1jhnPGjf6
FYzt07265s2NK0RyZ8ZxuPwjl5+wPF4RGwawSHG6U01AiEPqqdB/u0Oht0Y37pgurd6wfC2oA210
bpja6XpF8VZLYsbBIOWfh8t138YTAJk8qS95obkV3nURHtBUHEDhxy5o+49QDNDDpqhbJgebJPbQ
RZpe/DLukOeEypL0ah/MQ6SxtqjkSzwcAEAm0+FXpt03JCTl1m55woU/pxvq3ITFOoPpHH2VCO9I
kzTi2lqy21fwSEbGCcz6zNLf1+/dTvr8EQByMeHTtPfFTa/WntOc148k3iaWVmqz+Uh+f5cGZq32
xcFtFGYmXrYVuENCF0W2TKuo8jJDjkrft0jeEDxV9A7BXK2Kl+9rBgDOrbbd9coyqwT2noUoHGuc
NQo1wrwtZCS6FmEhjZ2maaPTJDObS9DcUHzTaC1+hxJSyEbhpnNZ09Uxr4mTkbbpmqBSc+hWPD2p
MSVrEGtCH8PHhrE0FPvczGLlC1yoLyYVpmb8571Sc5b7aXOvZA+ifT+p/SmEu0sxanVW66oven0G
c88ZpRik5fQV22BZZrSNjauP7R85DrN2RIeqkEEsbyLRVfWF6yfq7RWHB0hCU1yGZEX05wTln5/i
5h30MwMAa1F3j5ES+/W/KdBuMz6kgG05KQCOWEoKniUDwrdiK3CPckXFSeR6h50M52XwE2LBf1dW
VBqXNrED6SJ8iVrKYlRfEUNsAWRaO10YK/AEPUR3VRlxkkiD0FvAMrLTl0R26pN5KKIXntQDnmnb
STbwkMnKMFymJfSPluH8xOkh8FdOCsbVldxogBXB4e0XVzicuDyZuhvkcEZUx6501m5jR3dt+vLG
a0VeurBEvbI6J7iAkxGtYEV1qttWbwhkpRwd2vwmxTLC92ZpLPHUE5SPR2MVh1ZJVcNeExLcj1kR
MFbKV2I3dY9Lp1ko6Kn7xonW/a89gkGvX7FqTC5SJHNTWJ0lW7BOTQaD/FN+cH0HStW4iEEKrzPJ
eEdm3bw8gJxc0lBTYyOamxOfT84M5un2RaKow0GxYAn3JohL7GaH1iHgHC8npnyIljkkP8P1Uvev
doGQDv2dOVb5CAJm8dzcw6Q4A8j1AnQDCyhBW9+JsIOS3OYiMR4xR1wgLBhxOOoqXVFN4k3/11pc
31c7y92FWZQnT+uinYd9Owaj5se6tzSEwaUtuIX88goR3STPFECN/b2FslDTU5tb6f+j+VwNcxyf
pamsB5CBWksXVSAhTDcPiaHtOxBh2sytloud7Dr9Ht5MmCIISaPSalH4vOZ/N/NGmzptVdGSk18C
1yJVUHcjzO+tzWbbvlzxdXQ9tZUuwvciVF+65eWt8RyGNFxSooThoeQNO75KQwY5rSBF71MyinAA
ivOfErCw3DilROn2ur5PoiPSc+g5zLHx0oIhX8MgIPTcPTi1ExihP22Df6e1W1E2Cq/D/hhNdiQU
YVMWwQxEYEunUSfY/aiZOgHqfTpZfXPydN1AECtlErWX5VAr78DekBluMIysNSSlt8uNqjJWqS1T
9BOtXEuJLvnbq8CUvfyS8llYumTvGphAyCp8Hi09vG6gxFiPqLhG56wMGOmu3A2LMfqJxpcOPQ98
bpNZoCdHvmZ7+Q4OQUPy2WLq8hRjSCZx64yTgMB/v73lGo5g0Em9+/Lg4Myexai2DXDVrxQpH71l
Jk4qOTwARDGl6QXZ9JlXUaOZaEDI1VC+dDYaxruI/OradATZdqevf2ySgZcWYQXlTrd3N8MwHS3Q
MCsRQ5aEF9S7/eoGL9t1vdfqK6kCXEiCV/tKpDZwEZFDyglGWT3pohWS7gT4y6jjy0G4/HPlh6E+
ZpGo7xfa9PiSzBTB2nDotudJDJRBi1N15PDXHHRqrLYjeIcyxZFyFGFSraW/qKW6r+5h4ZmfYtVE
zWicVg2uGfAvzFLU/HqDamsKbazALxPt/weJjn6+z05MuDBUfcVqQCRbSI5bAsJsWawru6TFp/b9
pdqEarjOICeu0FxRC99B7LL3NK7uVRITHhxCTHiLdW/hrw+3vJ+xOyoowhCkFkl5NtDvQdVmqc/i
eM1Vbh7qktz1qqVx1rWslLgTFYCpm+uoLfMAGCHf/9ZZS0SUimGPb4YqFr/a9TuriJNx2yGf1AqH
tUuJ7KDf/zE6DbR+wydBJloA1beUI6ZXgDNpqk8gt8w6PikB4ypt61nnyNQ3lw9SymF+RcGtj6mQ
KxmK0lJ8lo4TugwTqVyVWz8E8z3pCB1ZrJgi42bUs43OO79FrzLOijVso95m/aR1egQ7Xl2o5xwh
ib21g1LJLdfvFbYXaQN+7qxB0AMDl/EuUYHtnbd3QuMkyxTJpqoTuXPjIOj6Fz/fiv9Jc2QdC/WM
8dBsFvI1Cwg3CZs5HI6BbyYP4qCCdIcLkk/nKp6bHJ/mF+TpaAWdkbF6DJXFGFIYoYaMNREl976p
pk9marEUQl8qi8JivIMVPvwR8RQVZrOPILu+gRNjJys9uoQ35i/wngWpREIRbOAeoSGc5KwIgbnB
Hs+2kA0gW4AfqOOsdztm8tPvfATeIw8/xBoditgc3b7V7lAkZvz9nKppT4OMSoLek7D31pzQk4BK
WaKjQ3JI0tjW0NaQ7hf2829BW8H3EnWFX2sA28mtLtOYEZ6trNZ/hsc/uj0cYVKHL3X7JC8/FC4i
NRsCoE+TM2g3DteQiIRm6mqFc+TxCvbeDsBDWT4kcNRiKQRxjOZeJISJSBKS1EVf1B+nLugbUbiQ
68v0ywyL/Vvz11bo/IIKyDoApPQlV55hqv3CF5BU48bZgUVsexsqOfPRMsG3v0w9gCf7+6lPrUbB
uHJrjjfATSuaUmJT81VQP2RHRZkWNSMoIxSyUbHuxOCqngIe13whHQkAY4DxJ/+oCmfvv07KqTzE
OAON+DbeG7Dyf6rx3THKClbg6oYYhLXySK6pm6JOsUpB49wzB710LdjOfUAJ4w1xwRGOb18Ks143
C5+DseNAlzqgmEdjh+GqHaLIvEbGrJhOaamvHMcCouFrwg22xilyxDolN+VMHEKEYHwzGDQbkJKo
V5czIRQFVgJB9zNDfBeZPEy8Dh8EFrrzggyRN1YnAuk+vI3oZFxQHvf8X3mLaUSU8W6EcyuCwGdN
g3uqjXwEDoCodTgSHGUnyxXriZdA8OToYAFkWkCia7KWDP5wwNJQkNXvdz7rA0M9d9cL0peLz/XW
zn1cB7LtPH+GtdidRJKukd2te7HrNT7DdGf2e7sSBl/cbswYjLCjt0iqQWhG6XEdHVUPkXWz5qUX
S75PQx+K/N5mqkfK3na0iuXqdQpEbMs5f5H/9io9WXBYiT9st896dwSoxUSaxjPWjTSm3iq/WBni
X3DyzG7nkhPMeQxA4ZrgVVDDF6HfQAY5QuHpkqC3+2tiZPDszn6f9v8rJrkG9FwO4nPlZ9EjAk3c
La/cD4PcDsLNV7oSxLNg26fADxWZn7xHoa+X48o46RnLD3I7GrnIi7papNV8LhaR0xlUpqGhT7Sx
vd++kWOzt3feJuDZnNLD3hjLepl+1QZ1fdi2UJQtVGWw6tgNRsKHl77XdLp6KFYdJl2mKwlSB9IX
yJFFbxHHtSQ40IDFub657ETx4OX0kQDCfeuXY/AfSpvyoJOy+aes0AG6SkeFaUG+WZLpV3j9W3Dt
q5wuU/HsjbCyh19Z3C2RF5xAWK7W4LTSgoH/Z/ApzGLi+PReFP15WfoAzI4hvZ3q4GI3sStAIWWk
d4jPztQXblKKQBxsSkxesYbH01iQrXkRB3w5HNmrNE/xC/uLextLvWw27i0ELKVZyCl51TRu5HmS
VfKYsTIYw2tep2X1exy95yTIZwSdXA6gz9MLEIM3ZLtMz5dJQnOkVa5KpkvO5qEgMblKN7NplJIq
nVgtZxhFGcyEn9wgAUJ/iYmWIN3AGhFE3/V8UnW4wmhNccEioXAcgU4Ngf9BC/lZrLxs9XFY9UpX
oFrsEHxGM9WlvmgppX9GGBSTS+bJ1GJpeGBuCeFY5Z+OlhQ2xpcHlE2imWal54bfRKvCVcE9ZwX0
EmUsr45affojhByIyBgvzpwjuSx53YOzu1AOJqmhVycqOD8D7KKwrAKiPEjI0ognZvDLUIGqUF6W
A2mLMPJTmUZ1NBrVp6RHMK+iXG4htWu4U5HgCiupdTB1JQWr082kKlQYPwjFoWk9HONXg2wzlnWO
cbY511AhFQVZYl2DoY+REeqg0UmVfmzF6c/8ioSlPjCem4+37De7MtIgNJK5038cqW5QSpOhq9p0
zUXxlXMvyt4Rra7Mr742+aJeNjxtk+cbQ+sWi+En32s7VY3K4YTW6gYjLZmBJPppXO6k3zg/F8iM
xlN2rWiVSZXV8d5Ivh26903uCz290BeUz93BHC6ZS6HYPFKUfoZeXgFy6f8K2uyS+BFXSjZrNGHZ
HLIZK2J99WAziiYVGJquqAtiXDKdWFzNhc6trjnQlGXFZL7eSflQNjs2WdwOzerXhcWay1SkEX2G
iDTmwtz+0I3nOPP54pEjH64jwc0J2T4Z2mwBSGMz0ilFZ79lLPWS4nn7tmVk7jBaQzC9p5H4/s8z
6rodwp9zxRYnUe+FosRLHnSTNplw3fBA+r0IWmAUqlzKeczm+jaSJEYIjFHPzo/+38o2U72eJLsC
tfTsBcbI4VNrr/W2Cn9c5hXAUg0LQwmXxv6HNv7YCNfXguTem4eYyipEj0Srm1XPuWlhWZhgzP00
7qLkzJxdUZ2A3F7eSdUSfw7j4DUdDTsgkVcwthqPJbnqDpEpGNFpkZvBF+USIZDZf96RE5QZGonV
vJP4p9HgOXH0OD+fLIZRoLhcby6IiJm+AS2BbBiiwKN9LdqNS0FOzeTgaXhJ+rT+HjOctohY2Zqo
/ld6UqJ5yR7Us3Tixwk9dEfgTl6WlyhdAHp+87FBM1uMkIGLS5ukwS8REwR5/vlEyRLH5tTCZLRL
kF43pc5b6CyvbFYDjs3yg3zzjBCX32ldJTUKn+BxvYlMjIVbv6HKVXQqwsR75x+1NGwKblX9tiAX
sgtn73N2RaizTj4UJu5GM+sSVU78JzWDMriJu46lk/nzGBigkDyCWcknJEkqbPphdSJVqJ+RitJ+
iP3ezSLJagbB9WZvAEcoKECj/2Jg5WKb/PmFUVHziKnjPgnxTqXItY99BhPDw8QT7yFW5Y4IIzB1
Gc4k9ZfLmopMOENz5MA23Zc8RLFUlG3p7dTuQaf9I1XTTI+/8qzWB1Wj3COkW1fF9Eq0UH3ARgRa
sm5XiVMMx4grJOP8OLobpMqAl6Jy4sm7X+lFkPqYJQvac0f7RN+DHMDYtIkgCNRFAyJhu1YSljaH
n6ydkuLlaQ+un6SFj+4kTJXXOZLsVFoWHb5acjI7QudSpaJDjdF+0k/Jy3wugym4pZQfOCW1yypf
0fZJfXfJlWOzdpgDmBkkkzPuCM4HuJ4/IgAHuFtMNTERzBk1sTnseqM9Bli0hy2C3nZypqoMC19D
0/VCehfPBVG3P/ZWmycXhVv7cno7G5uf8SMFWzjdNXlTkHoBKqEryjfhUaLaMrqzluAmHewCp0oT
5dqza9971rd2WKA3drSuQM71iTPESQq/oQxmHgtgzs3jArHKIMXjayVPRnkjydjewXF+bZgjZ1an
B1JOpXK75fQ4EkfJPpxhZ60jqKUx0NT2tOb62Gf9bluOQcdpBO5Xlj1vi4Jm4K44ITEjVAfQL9MU
p+fNZgkESdREx4W44kUR6echpQtN5HPmRq3UHBU4uPjNNS7MVxhiHGxq7DPVnvVjyp30J1sXV4QG
oBnMZv8GRUgHP9HBvngZYCDqecYG+mtyzkZSTlxbOWabs+Vjbcer2XjxcxIDjQ5GmLmWnTy3LEji
PTeeE+kaKYTPsKwtzpELaRQBAd3/nqGM2iCpMObpkQATVJUZY3lVbbQyHA4ZgsSCOEVA7VZAdRt8
uxxMvqtUyDnpHBJFgm07haj6WErFDA/q71GQFKl7tYA5p7J0JzQYAEm2BYII64sUqpnM3tks2lcs
J91hR6ZGppD0j5/Q7Ldx+Zs0gh+G+d/DEKizA6s/MAuhUiIZd0Y098anlbEDq2sAcC7fTUlCc9nh
d/xbPXtSfpsgxA1EMeFwy/SJpLw1YzaaGoj51yPeJYX+ueuXG+ti9+THqpvxQadS8y2CYj2mRxd7
YRBpQLLmX+CavmM4JMxs9tjXiHfPp0/D+gRTL8/tLbxug7bduhnImAA2eORmatFKuBZhFCxzt1Ye
/65AM4/e0xBPyUn83Pzr6JO3Gs+/gzFcbEHThAhlhTqV+MiMWhj2tbfakxJw1z+Q5A5LrwRglO4I
hjRkSI7TrX+3xW30QY4wRbDYR/XBmQOiz4ithG51WDko88ntdUCP+CU4GtLtCKN+cnq+Lt7W7FPE
0fd473pI2jg6d11o2ar9Ahhv6NKdF6gMqpqiv7zqg3rl5ZBB0Hg1CFrmWRXePL1dIc4X0RIWT05k
Lx04kZyjTXUaJsBaCYbSu1CJBpbM7RuHSsb35/tVC/t0XoyoRGLh3hIrY+dgftTIrgveWCgvJRJL
3p0iG+1xK74SkrrpX2g4jPOIizjyQtc7jHD52y3CNZQSuQ4zIiK6DZ6002u1fNOP3sC3F2wO/E/K
cm7n5YyisikBKNf3a80oNURq7TLUoiVx4/hFaVY5+vHA+8xnISkvy0hW4TPnoxosjJ5BnJsfIhuP
mafo3Q3sNyW/7g0jvhcyehaZe8WQf7KLychGgmsoFV/DmWcdsKB3xhY7sUI1zPPu5qE3cI3/OKGD
1O3kYsnNjs1jMsy/HBRXqyLXJzbOe++jWfo9guEv5tku7sd13UQCBSQxeVJo4phPM4qOzq3mnG3x
4TQvAoF8J68z+qn3H/AR3javP1KKeoD8EQWZYjZMHiy1SRNmcU67eIFpA92a+bYnzRppxZciIDPA
JXdnhrxSQuivCjGdyrJDAhIyWbd1v0UTFzrN5TqcD0ea1VryKJxIjdqHQGU+Ipkau2hE1Mvb9aBg
k4aa/wVwrCQ9IE+AHTGrUfZAD8lWzG+jmJ7RMRv/L0GBV1Sea4uA0KOsdD9+6mOpcJfNv0huAOIU
NnNvAQvO/22uILzC3xxlE4GGutzR3bnlOwq3Qjm0DACIqt5AS8qJl0L1HrUQcprP+2prrDsQufn4
deMkFUSwad03F4FJIPhtfVhWcT9pMD90Goq49/6A4O7QePP+IZIvUr5qgV/O8adym4td/EOt6zgV
r/rXUeokMt0qylD79YrdpAwB0W+Z1kNY3LKkr6XXm2EcBoZ+I+1+hiEWtJI54xoGg5XTntFOpMo/
25xSS7zcBFpyK1PAU+oEr3zEVCqzEqxbbXPzcAvOQbFaUJpQjKK/hygmkY4r6G84lqA/oMpwtPIZ
wLdARLKlkTMByb8vdkWtORy1gW8sjf10dH52cLxN78sRMsQy9MrZVzwO3kN/TpuNd7XRlPss8+wV
a17fIRhfO0gQ/q3r53xF2lil8r1M0iwqS2GOzYBS2OOmm1ggX7nNJuXJy0dL8FLKLmpzW9199z//
hTKj2dQNS1Kp4TJqNRiyx2Jrj80iGmtSiIzNVqOHfArbEX4lU1IqlB690JA/8okEYNFjF80uJ2fu
hR+qE9yixmRwwYHvrXMYygg6fIKofGdQAEA340o3psixxl508gyP/Wj+Krvso+mLzXWogcg1K+Hw
Z39RI9TXpQ1kVw+QKNhCsxPA7naU21qvbLezDuWGP3g+4HRGiGZ+VdwMSLSVqRws1s7Fqlx/8RUo
O/m3oxh2deGksFODz0Qv9jM2jZNIn0P4+ji6LrR4Ohx2QcBjNZbqMnISOEQ1RkvABllGEw+ULnSV
AiKiMZLGqUD9vk3o/Qu+1fzujba8xs7674sdUP8vMpuaFkYI/oXE2bqF4QBks84RbvZzBXePEYul
34fAzCLEOlGLey+TN6HsJyQk6KGl/C3SAXOHUpM0IwUr9k7f80WU7f4cFM+XB8JP20aHn986RVtJ
uRqfXSQppVSLrEA7y4urSJuJcX0s6l+lxIjfkpGYedvLZcvOH/DkDAs+oDUmwhjSckT1y1XPa9zj
90uXBH85OOnOAirADk+/kVrmfK+UqjSbf5Pt0CL4QjONEggIFMuV340mvOpt38V0wNORZyBCFANg
DZ4gT+opfJCtycWQwfpfdhEHPx8K8w77yJg/PiPJxbcL95odAT9jiGGUILWHetjYUD6O+5NPZFuc
4NLI18Md1vjqJwQFa1nKFMzMowVS10eit7GvsYz4lckPGVm6OkwSkTySoWnhv+Cw/rcF7TCT6+0o
zKIatWQFLdazzxCVLHHT+UQSKzx5+AkCGtDpM4gXC+YzR2w2JCeFt17S+U/N3vlRVYuzAMLD8U8p
KipwZpo53UyS8T0pfL3P0VYEai5Dqc6VUV0FXCI7fcdPjvfBZ4sAev/S4mxQZLlM1sArv2pt/ReS
N7+VVKGJjYWHlUaH4debEgMJDiiyD0GRUtnWZIL0hWvxS+L1BDAS/oSsmXC/FSi0T47WdxqEzg9S
Nfw9wXNnKM3K7YFyH2EOVzajznRzel1XrviBGPupKtEh4lYV5SrVyKkam9lnBrOLErSoPc6ISVFG
0ulyxyX7hgG0D4V02psDJmswz3Vxyq/Bv+vZj85n98Dvo/ydaqf7omTqXdZrRSWN87BAGoOGsYaS
S+0ZMrDwHgHImm2+PIlnajPZPAf6bSk/Ga4UPfvKbwf/l1nuPNT18LJclkxNEeKYcfV0TEqHXFVk
Y23Uj6qNfp7kMwD3Z2U4FEX3pBvm2JBxendoo288g/oLn7Vs8sU8BqsBxDOBpsYCy+ktT1t4cRJ4
IAf8xj7cfV7uIR2C4NUMyIdI++xEww6AvtE2Rh7OBLBNbaN8pIIKVPTza5pNNqb7bXqfSEPk9nKx
Bt1yhqCEAiOWhfayoZL+scYPfWM/V7AgbSnPOSUYIUIjBu2IJHmyXGY5FqB+Lmkaovo/OQ998KwM
fUqhtGELjx1jhbVOG8e9p6b1DyHDHYpbZNGfM5/EUoss5ik+G+5gAfH+RxuseB/18ZtHrBTtEnUq
VkVJUrRXRBGVsZuBvTHwvmeYTD0p45qIFQFw76Po2Xdnrt6k1oFL9y9qPGpldmBw/o9feCGvCnfz
h8J25FssJWObTC7MjQxM9q1NDgxs0lPDRWCxtSWAiDdVPAv0Zv6pSs6EtaYq9FL7+XM0nef1wYCn
fzCOM28KkkLKTFBCyymVphNlASPWBcHsHYhqzX1/sHi30qoiOkrJ2NY2U/8dhzdUUAhK3PfHllKc
q3/1yPFrKg6qvkCZnZl3xbQSppVFwLJ7ZVYTVY/jLC/a050UWvpZNqaNQieXJWpd7KAA8g1m0Ej3
gWSxLY0Vuy3ymw6OctRaqlzejd3RC9mAajF5/OMuggDtGGb1HUJ5yZ3PhfBQvhTYjf5p9/j5yM60
0BOOB1YwOghQB50R3d7yDix+PDOl/OklbtJ7AiMGJvZMIqmMX+EFzRJMajifqENvwBho6yExXHAy
gIzWo7r/mJXiMiVjaJLF2GMT3uxxrjhamoiCSo6rkE4NKV+HFyZWH/qegogeOvB/hsXYLbgwh4P2
MhIwFCxaCboALFhzR+z4iJhu/F9spqzxSXfZijiJkpgE+v70EnOZ6xbQCCl5DI1+HUABFR7o6KFZ
rXNuSudrprG/4IAsRZUDn7Cn7KQRr2I4YWXV4rKEeJ/RF5Wf8aWkMCuQ+biixi4hRtWNcfZu8C0I
kSTUPe5uJoOe37kHxaKSpok8cyCVh2N6/egXuyVU9RnTcG1jnYXNVY2deqnYcJRAUG60LAcyJTWr
QaHU6+/WCq1xn8UErzcUgDF/FfhmNo5ctmc2QhlWP1Fv3AnIN77gFu0CmffpTd5FYQe5nLO6M2lu
rhmnigCf2VL4iiLyi/bRqdDXrA+3mOVoZIYsZ7bB+Nkpj+TtWX2e1rVIkkz4JW5hxW29XmNrIWlv
s5cIfsrXvSvY+pbteKNIAo2mWey/5/HVUOUVm4HQLEp2bqTG1c7mCkcn1dSVqGF+etq+Lj22ZJsf
CsYnXib4BAQCEkgnHwCWO0dCC7KXl8wz0/34bV6XJ5mSn4BdG6Z3VobZIY1Y3e9ln6+kHrMi8IB7
8Ad+l4zFik+2mpyA+CVJQihfyCwW5LJmbiaO/9HS9j60chjsipVuJjZQHKowUeRP8FzbqZxoeUYw
NIOcDRLbtGTyneCi2OlXnQeCuHU+NYGBd07ObNmStXXx5Se2yILWLXA70OuLxWkKTsV7BPMb8iWe
KvIow06hRjWnmqLcNbzxBQeZu4o2TDwlJVJHTRZJlnXaTkCBKNGA8CHzU+6Zznx2SUu/0X0FOm8U
vzyhPtgo/G8qi/B0nmBqYczjO0bDqu+EB4Nth9ZtkA1+UbFKJtJ/sE+eSRWogjzr7ekF0Zylxr0+
5LCAs4uxcxrhS7dGNGTI
`protect end_protected
