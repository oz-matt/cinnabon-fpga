-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
iJFUnbcagrWGTV6qzhve3XaTBUx12hXh1FPih86v10tgdeBYkRzAWqcNingAlKxlycnj5Mj9l5WV
+8ObbOfthYZAQDEuknzVUR6PDdTImhQDPDqdSH9HJ6/9KsGV4yu4GmEmzja+9ZAkjDzFMwUh9nXb
Rn1hieYgVcyzD5KsrYeODoZSv0m0o9lnV7JbCQkyVdxAq9P1Eru3Lur19qlEFv7rcDihgSGday0M
RVw0hY63KzG92yvOfXRHVQ/voUPD8XxZ4cf5wmY2080c5XwWOWkm78kFYuoggUsu5ImXrlMk2n5F
YSi69XZrZdBRuryQi8asC5mi2z4omJ/bZrzc8Q==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 45120)
`protect data_block
AXPiotDfiTTLOR0MqnD27KdgGgsj16aMplnr9plBx1nV8DojtnJMdfzH2Vt0ONZpjbje6VChnVqY
PsXC10nCzjXGkfRZESO73pOlAaDYtApXZMKHIlhBQ88BX1Qf/2SkkwCVWi36+DHk5Ov7TdmFALuX
dK+88RE4L0ko/e8BIQhTJHfqN3JYblbZJF71MTWKedFJ42rwBz1XDFI9n/ppMcYwe14SJfpzKoMI
OvfZOCJ+J7Xz+RJUveKgOF9+Sd/NwJYIP7AkJzhhRyR2xNS0cJ3HK1VS1nROJ5jjRTnwWhVt5a+W
8d0d2iG+sJFR4g0fwA/dLomrmml4xSAEVx9n9UKtfA2UdD0do2Y1iixwO2r91HJqQA0yXeRglrlb
WNCQpCipB7hQYKa2C3Hhcx2VayIGWpVy1GRAOKb14fHF5wtNsCV/3E1QDvutQSihUO2hRUZipPqL
VEqY6Oc5ARodN56o/hgSguTwVRCh+XcR4UiKOslH3HRrqowjzI4BLqEEV0y04TGkWdFHcKYq/Izm
p63pzmhjs2nu4BUs9Gvnbgd5HauvwdGTWU791xMdq0MK0zwe47SxQjcQNLQrXgupFodCX2CPGSDN
S66APD7SxBBaepH3CFxxbhjNzE6RiElrE5u+Mnt8cK5QvAlzqTbNXNq2xQWvY9wupdq6WFEu7pbD
yqTODFSt1vmgVxt5Jw9+otZp/2TO/9hO1v5Nge0JjTOwmylgghMGi+A3J/t8mFCfKOgHNjPDfTLp
O8RgU8DGL/4OR65jo4xWLLY7AJa4PCZSzs/G1rOgCZb38Ho4/uhlFyYpJJ0rxTf+nQdjwbhUscHB
BnHh+zDqCFjCkYp6UhJa5Pv9mp3qH5F4tIKUGi0r9Xeb5QEnykMilbVTW7tIpZLo7wVLb3/AZi79
XVRVRc6QJg64NmbVgrGtO5sWoE55eg4RXTS6tqVPxMJO48UlqkuBT7OfU+WVDMiPufVOqxNi4Tia
Ngcx3uGZ5OP/RzBide+P/6VCh2BZ6SZuOCD5nk2Y0SlAWOA+LW3qO98jdSyu4M1hA/BBp+CSTKc4
7szhN52AVaYuA2P3eRX5RZyNBjC/MkvlFnWMDbb3JF6Ea39PTbTHHV01b28v6OHg9fZ5SLsekKqs
5jqLhTKHiMEpZUX8trtQfSnLvqJTdENCS3a0KPrSoHpJWddgeeE3/q6ldEKlgUV/OpIjyjt8x17h
GuU6nQUkKqz9VGXiPM9UlmkOkb1e94AjlMU4zH27OsA9cnx4veODBGlVN5x/nlW4prdUh79SPR88
2HalmjgUz8NCKj0ilmPp/QUotLdBm2txEwO5TBsxvGtayPiCiIbC0AEPKuOp8YS1dK8VS02I/ADM
/DCIDTryUJmrN+CFrUbRn82/+kjlABFsTfwgWL+CbwO5zHl7IxjtwwKp5omozazClS7cZlLIyazY
NjgzCbhRf3ThkzeKmGq50N4+VRFD7Jddj++ni/yGUHb42DvlUV2Lm4mvXIZ1qcJwjX/9GxjRBkss
Z5uHJ2kN18bskgZPJDOr5WDZJBzdjoPHmZfwKCFZtT8HChFpBH/IBU2KwkfJF/K8rd1Af7aWRXwR
OP5xIOQS/msDvv8Rt1KNOTSB93w02Z7OchxtX4XAxNsRcjiSmH+rD3WvbGLlugs5Vxq8gR7Vixnq
c9vO84aIAw0+Y5RiA99Rj20HhumRLwYUyu4M0c+tJ2ALe39u/5d3AUODrd+XbV97lUv8pEFz8Inm
CPskxf/u2ZAQTOL0De2PRV6OQAjPmlQTY/VGYYuH9koouFFNXPVex/RqR3PHHoJSs15HJCqqrdLg
sCFZYqpyG6fDcKCA+9dQ9JUt9YpuB2Zn4ZrMHMb0w2CgTNlaMsDI1h4wKcOHwJ7vgR3L9XksmhMr
6eCZnY7kDW3I/ZsRONFj7N31LWBhY4jJmQuNvIaqj6S0qgDaX7o0sH8+TmeCZQuG9trePIsaMfjt
ud0Uf9ZxLBaENSHMbhP9+XyCcWA0NCtRMuCPGlhkCJZYteeXCpI3tF8bLnH7JABrwO5ZYafjkdby
KAh8NMOtfaMtbQV9+IgLNWBtFdGBiJYEOO05wZGV2oXsyaS87BDmFmLtivZ3qg9dB76/njrHgJ6S
GH4fH+r3rphVEjM1WkYjGGh0PI1/h3UDTiPpN99k8KPXwdmyPmumCteRfYibeUGyDEov4KGwitZz
z6N3Op09e72H18ZoTNfzfujbdnOM907cnVVxfMZvtNGJIZeL6a7YDiPHJjLjI72kPjplC+drc3eB
tD0eeBsQC4SXufEqkhie296ObN6O+G+glBCBTAB0Cdq9khx9nChC7eVkkaaC7I5hph738OYmP5kp
koIydFfl1tKfHfJXMN03xFDl38qgYvGE6V2hT8UqwhVRXJ9FtbX+mqPzOEv4UnJypNEn/kWcTCIp
WJrJiKVSJeAWJMhRYu9AW6W/bGeIZ1x6N/J6/lMLIpk/y39+NQVUByxfZ95Ea1+GFahCT/jMMBSk
REjdW9cOBicb32lO/kea1lridZZcvNsr5XPwPRJtklYmo4ynzXWtR8pb/uxM+kxTosa5tG8TpaY5
n63hcJYh1jklMNB9ctvAhPcgvjMYPlzk7Asi1eBj4B7wVOHeePARhTd6LLLl8p4pR26Q4CHyx4pq
nGsagaH5sslu/ABTAu3LkbZu+zSGmv37B8gILrBQADMeeTXk0v6lDhOeSqguyPzKt6kRDHrwDTCK
GkZm054UlQ7vTTU2BFxVZkzBSHtSsHriocwTpgGvilrd1ioWYi/o93u63WR9YznsSzspay/I3D0I
HtvORllBbiohvesFt+bZWD58yMZrr9qIXBv61XYtZPTmadRInBuWSuDNPe+DI7OCxxYkS3NUD5Qq
fqQuuzyhhXEZ+7S7DaANhbQEFEhu1iu03+JU96LNA7+ntwmaGb2KjCdwXq4DPboxiTZkeyUofs0t
UwcbOv/YgDzD+kkTrxUmphZweuyiXVioqwN8mxtpkOOptN8G+lJRj6Y+xC8c/6fYQPCWI3nUsG0U
PUh2yrNusa3V8JICvWXC32utj2+GLdmI6r/hlURVKO+rssNhCQvfiBGBK5RWGDvRjYRHYws+eCsD
l0eNhQ9aFmyzTBZlavOFiPtaO6z5Of7rGsb/dCkbFcfMMM6pfjTG21KKkSkScEv9XmWM53uM7wpS
cR6ImV38EYPz3mLUVmuDrLX5bcGMNYk07PtCHY5SNkJrLxlKG5d5Yj28THF/THE9YI3OsFBptmQu
4fB7u2vSvJ6Vrc1Pnnr+4IVFFdDkTM8f7IHnRpaiZAznnko/1v7sg5JirEcnSEAZS4znuO2+3eR8
hAqCnqJw7svIVZHc26N0UPPC62oCLFXOL0PK6ZzCFbm1BbeUanma1288WhUlLYtMp79x4qPmD7M1
zTb3MWS2aAbgaKz+xWlqwJY77YBo3z1RWa+PgjwygDiZOnruc8h3q7VsJ7H7EvYJg+TPe5RJTQns
CkZDp4G3JH/7Y2wPSc2U2b+F4YztqaZmDkrxrcIhvlcf6Z3yFtg211WOlrbT3JTt8rctYCKpx+u5
Ug1Vt9PgN+JzXkUci1F2YRhNnwBM8PHlECMkB+2dWOo4PrPxV6XQzFS/YRfP65gxJ4qhb6wJycIa
KzVFjvS7aVbidAU7Md+euC5DqN4et/gxsg6Ey+1ewvCVnEuTdT6imBuXcefxzVPI1TZTdxRWDzGj
xzwwXwUXo+FX3P2Is1MUgW6/nfoI0djU4Y0V6ZoKxD7ZNIo662qmRXLvac+6mck7DHuwdVeX1Ky1
iN47YpPQsGfZEwoIi4wZNrTfTiUrvvSHjKauskj/LUDf3hKV0/floCxaa0fMARm8OMOZcYt+16fG
L/PpglaUV5/QYvKbI+ICahmYEHCPRqdkQ7+CgpXAWfn/ik6p+M7E/1PBuHxKPEiSS3xn2l5/U5s7
PGh46UF4/LmtxJlH8G6GXl088+t+iqnRAOrR8OJ2mFLcixrrFPBxiuSX5vif56TWnYKxnpDrDTF7
CfZqD/+Hq//Qbflqvt5vwsaZxvHi00BvzdMKwvFfK+gV0fukkbqKsigKYXAR6lUNEmcJT12ZQ+KD
JCHYHSsat9jNzTi147my490dBHHQVp8VFwS2DE03w/DPrSbLSRd2X9OOmvSscnT3YMGPVPLmVGJU
TQaDRqRVFhqO/0hExANufuM3l/V6a6LVG8VqSysSixlsaGHmybBJzi9w63QA8kNQAkcM8Roa1uPM
bmz6nYnv0+dxYe0KzoulF8D9ZSL7VWPqutP3n5+7bJxfR+HLiCtp+ghs6vLmc1/pS3JjrO8O4sp9
jKtQfkvld9vZqdDiLuJfFy3ZkHXtb2ccXxR7y7xOoHZYuVpnbG+mzLp+mscqkYenWNkY4UOP9/sx
K19C2bkfldg4hk3DIVyhryBpaaNiA/U8RHzcwXHEVAES++ytSnB5wNCZxMxRdxl3zgoWt35BD200
j+ttXftLYQn8vLm3+mAYkbPXch1an7ZAud6SsMM5q3zJ/84hao5WPAhti7+G4n2p8X5H4MOJNQZ4
bszDS3q4VlH5YrSG8Lbn3D/opZ6cZufc+7xf9sAJYtqj8TJ9is/j+1AkVAQQGvyN+z3LGvx8N72b
7mapkE1Yi2f+X1oX8Ftpk8K6CWR0WE4PyglyXNX1Gj1Iv4PnW6A3uYLCZPcBfYhguntwvvEBx+by
DCL2z8jsxpVaW9PHkYF91SyHbe9fyvKB9RRh4vLrPXDd8cj3NSGW5IJQZFiW5k9NbdRdvrnFFDB9
BbMg09H2+02jchPiDaD6L52A1u+l3ndJ6oEJwVgjNl5djRayPsfz65BSr9sRcW8lIRhzGlFqxMAu
XmWX2k5J68+9zfLq+kqEOeSikZ09MGkCVbjoA+3CfhGu4JNofw1FKSOQ3CyXQG8oFJtRNvNJlpIz
Gle2BNYDsnlDNkQa+y+9wU+vlFoebVUxPxoqjNMXfNctOO8Cy5eqpk8mRuuViPVBCPtYzJYiEeBq
p8ejq8wcGyhXe7Al8IBkX1OUJSMTleBBJKIMRw0DPkLzX/qBVjQ6EgPKHb2d5gmp7gPAgGr8nPO6
VtWSr6N9udEpiW8ch1t7s+MVlr0Dt5xC/XOj+D7yHlJj94yHwACTddUhJfyz7v127CNWfFcAuhRs
+mvHlJGcX24hx9q6sBjOgvH5SzR2dLOgyujAnHt6HbKt3eY2+TFADz/4RR8k4tNQfDsRG55AP7cG
43I11VCKvAG9/Gm3NmjKa1Rx+n83+pgz7d/3f+pl8Cou+Vw66SlX807dI4gwfjs8PAHfk0lwAXIq
Z7rUomcpu2rlXFeAx1VmTg9XgADYEZHS6Xpnp5UXiZaESsFQ5m9XqZkBPDg8aHQOWdPdtMslnMYc
sfEUOAxEvNvVlys0vX9ul/y+TnLUyeouJnBB9smdt+b2HMOdOQPSXPOuQkjVp4Nu5DPwgpdQBCyk
CqKuA5xrxLm7OkrZbthx94yGXoPukH08lfQwiom4Xvuo/P/P0qkMtF38ImzEUiB9uQcQ102snbTC
iTb+NqjcRZRniWiodRsiufd+ZWtG3IeI/z/T2MusQL/3jtWQHRomQfvqcqL0YKr4kAqnPrvq6lE+
TCFrVoTAxxXYuY0BQrW8002i6wW0qd/7xWD2Bj9gzBdi1DdECk2pwWkdCec3tmF3WH3tD6Y38mDZ
vKVBpBnw2TgcnmmL9WgeMRi+w1+jYXy0UlyecV9MkrelSoLmocXb7CT0n9dHUg5Fo+PrhqEFMwPb
vPcdnvZRIWbP0gVglFOfgOIb1NojzWuYaOIdnbAyE23uHP9nTg9+acAf7kVTwUr29JXT9fVoH8OH
XW6slD0P/Ib0yDOwn4QFfzTXjTa2Os8dmcDB6/6DiCYlQ6vTQSbQB2gkaETiPtJvTMjlE//67NDq
NdFm2WzCMhKddD8z8sT7Gr3Q0l6a864Z/KYNXrLyB1FmGHXm/xQVJcHGu20kYDgFJqUPDeB9qNZd
sCZ8Sd/7OoPW8FGL5pmHyST8FUnPqLGkQxG6hp11JY+UJ0zpAjYqN4JmDivS6insnwPWpComn9/E
BBekIZBrastEm1zFF+HYDg5NF9+16mlOO2r7XHEqd/cMh3+XzwEkMMmF45/kQg+5Zp3TAJAV0MQY
ddDQA2no8Y2LZOGl5Nzslur4hIrRxSBh99t4jiEYhErP5hZp00OIMUXrFXlqUzIrgRBEsBEzYLfC
i0ifPBI+hQECKyxejZEhS4IvMJwshEkJCrF4KziDLhiGDSfoUHqoWdmX2ouqN4sWZZAEUS2c33uG
/D5x1MAe2rw1+iD0RiEKP6ebP5qg7MjxHehnAg851C5VHUBZweL4ylgBRmZHD+t/FVfmYH/w07gm
PS6cNGoHxD5dtFwoWE625eacFZyA0PeOBe5Vdcle1JvZsSO+8e6zBYweX7Ala+LufT529YAQ0LF+
jsbs701FZOgz2TGXMPjfZzbwD+iktMw8u6w/Y9/Ce9K7DfozZ7aOc3IxV+jKuSMUrj2eP1USq8cA
PfLEOIOkxY4mXEOnPPmN2cISyUvusol/+46uleqWwOTwQFqzT9gwJva1Zh7/0ZsRGEIEHeMIxjQj
0QCx+R9rF4sn3QVLDlfjeHgFR2gqZxAIBGA8hZqtbD9MLegLsvgTxmw5PLPqD7q6cyWdpqPhDidl
sqqaBb/Q/7JmDoZFrCMUmaMWFv0VecpWlnBOMeOeMXVQkznUTCogEEgNZT4RFt+IJPlK0UQvZLbq
6xDpyviqD0JSa6cKNifCqs42ETt6jXXHZOT/bWfO2neYObTfjpBYAwRQecUzYzm9rphceMmjw6SW
jfj065Eo2WGUZ1ZnUqPBpFcRrlEmZcOmUkt7KNAogwyNtCjJiYoaIyidVbZVPEt132q67uKqnTGo
a8kOQvo9wxO2NeNvaxSzDTOXFwZr0f4mGMl1xDlgohJVjjpsoLyawck28JnDTuGNQZy5vPCZk664
Xc4pc8S0Z5EKmmWeyZQQiuLTR9kb39hj93fNNK5czg0NgDsNNlNUeCyeNO4cijPmoLWScyffurh9
i+JzyLW6nJwRmMkF/5e4J0cGqxAgxpNq2d6hwBPPrVzBqpwtt0DP5ABkQhX7lZ19wg69lxKdC0ZJ
3MPlpIyblulMO67hfMQF9YWwy68krvRFHTYyZtPcPJQTpQ/eekVA3zbuS9+rvP4yXg8PrTcLZeH1
UUNOsUVDAiqXGOUM7UWbVlnW80LVjQ75ItdTy9fe2Je0PK6gi9JqHVJ0o+cypdY6DQwHeThvxWMs
qBbA3TeMX9qKyQsfE/bkWjex6wN7ugAPNpHCN2RYQt0ANAD3X/qGCP7NA3347BgNBVBewXUoBrrk
LTpeqg+iJuHTnsDCAxuxXbuac9othOiBXXPCc122SwE+M+EkPhde9a+kZtLof1x32fYb6Ro5cn1U
dWpZN8T2Noe3sEV5AiBOB7H7VGhkfpMR4f5Psh+rjEKeRQv13iP4nLrkaiAWipxM+E1qGGjgtV8N
MOeNWGe9OJdemaX9CXiALslsbBEhHfqHFWL7WK4ZREU9g1bXMO9A8k9BmRp53e1fIzLm9/yqXHd6
cU6ytih4gWyxg1feaPkadJEeO+MQpKNArbdxVVGFIrsGCgdrZCqREIY0x+Nn2SQkU/99zKZQNMmu
GZGcXudmZ47HCbLhywd2nTP/EC5Qi6jXhHsK1NjzAGefX+MPcm6Mex/P1hIY/L19sGnUFaM+W2Ek
dX1MtjgIPIl1GreY/N/3CA4oSlt/P2PbqWw/TmnS6o9D16mCAD/x/VKDyHumGY1QjzOq574hOUbV
qS5xPU58bZaRHxLXdHYgFgMTYKFPU9xYQM8Lasc7nrOEMgF3FGp1wkYh4vJwc0/kegSTVSSyBEhF
icBhJskf326Z361VkMgqWAG9r3bOafWQY0+Wm7/fFyJQ5QHF92/t4gfuA/bTwmxnTf3wdNXpubjg
YwLFrs9T29KwJ6ZqFfEoBp2+LFDogALBk91CoOHN36HW2kCn6lSqQkm5l5+JyQmNVd/AmzVz7omn
stmyeBdw2qF6KP0WAYNKLETexVlUgcZYFVocC5UORMvE9F+Ab56lvbm7utcNNVKkU9N8lE9lVAhr
AYUZczjaXPcZx8V418KVejFkQk4pA+Yxv2jJ4NzUkBs0gU+n3DdskoXdZyFXtLDJe2sFlF/7nLWi
nc/5RRix+IERPZ0FEaSiApyoq841TaARjIwcJmSVXFa0hXrPxJKX/QRCAmgjbKfeGz3Nz0yK6nm7
Zm6AZI+lgfrwPy9fTvCCf7eaEm9n1fTNMWF5KbZxTGapWzOwQNUhvUYhWTmKGpjvxY6hkFS047Lu
+b/dcVoGWB+cwRn6qbYZeVm9EGYIctz6FO3oXCqm7lIr0MWc1WJ/xXX9Snjhou3iUxb9PXmpH0QT
tM3Y/qENgJiyKoUQRk2ShLdb2qZXaOPuwIDfYuf/vJpXgEQUidjW4bxHjwa+6Nrxx2X1wYW/RKej
QpYmSHBflddJ2Boq7fPFW3aw0VYXems85NR55K3mdlJj0jTdYkvhTJY2Tv6JaouyID5sumkEzVDo
T0/c0ytx5E0djAanEULH3tEDc9RDlmynSs/WtiJwKEwVhlis24/uy/uLvHzZh1Nmtr8e+9jk6cw1
QnkigsSmXSGOFZjhe8/T/rAjItY5fANBS2Djk+YL0vcNDU5P6UXc4Fm2H563A/ZxUIr/2phE9LSm
FcPPPoKpP/3/UMBMwgQRVZjRCEGhBMamBcMqq2+HGopfszSgUb7X1QtuXkdXEDtNuOJ2wi+xfHdH
JR1FyXXQS0e+r/EsdbHX6Mj+N05c0+Y00Q1dZh4nQemLbJRAxlXRFpIJB6nzUVZ1UmnQgCwVUxWx
ugU2hh/jSkDYSEhZfj6QNQPB+cDE7W2mILq/Rsl64HXAgYohoJmkVlGL60Qb4xpnIzDu+I28zlhE
U0aw7bVPh/WGLmrSrz+0JRDS2bQBZHlYIxoDEWpiR4VBdqdYnWGhIKe2qkhU4mHQNnMMqDTvFvkJ
8ybOKFLfplq0tl+ARGumUFH6XEM7lCVBOV8HBv2Wy//9jSLWk0NslBGFMD3QleNsiOMionxzU7WC
PeGyM8mz4icCB/Ccj2j5d9wsNwf8RviFwe2AlHj6blixK8M0CV6rTjv5U4m9b3WcoNIaDormdIIh
mt8DIDcZrJ3ofRURYaoE8vyr912YwSPWtpfysvib9ZnEDjqQ41ujkCdnWsUR6N7ULx+A+UEvR2Ge
ctF1RdMzTyG618clfLS0gff7WfDSRAFnvorFIzl1bTAmeRKty0iMrE7SEMJQMw3LdgZfu/pGyujC
6XHyU/G8RxG6A2bLPlHDxGch2N485kgytZoN+tU7OMGMp2B2wKnLSs8zNiAka0/ttwJN0x+wHZHS
mqumjw9tMih08NgaPzBZ1RCQoXL7BKvsg92jtKImYSjCCcstfMqcrMmWbGgbGFchAsEJXB0pddTh
suLnIKGUigG7e2MNHY2bitYV3hs3W1ztKivYkTGNFV+iVC8z4xNwWIhgPDoWFtp4QXU5bS132rCj
Wee46MJ5LMsKq1r8tgBaGKbnjKhSasYFZ0t1xpCufipVFxMUueG4ZvqDeaebsAMNOCdc0XBQbWK2
eEBqIS7/Ou+fNtN7DNQ1N2+AyKu1yVh5PUAeLJsszm2ArAt2G03geQ1KYVnLWD1jyHek48MvnMaM
0/XNi/nYiuwOXcPzT31+uTW5VCC9X/QcDLbaI6enYLN4CCX+669MnVZFta+q49q0V23nXwsmhkr1
2cyrWAvWtuPM9foe3aUATBl16k4jvZwJ40qsyCp/AnMB3sZUtjjp20XHR/DklVfVWDW6Rcq0i9gO
JKnpwrXfLRt9a/6+Jay2kCsmxsVEoJSavCXR9TtVXv78q0wyXdI3Xi/qYQByNQLzInK74CxZsLjR
mEAEaeSxeIAUIlBc02ymOY/bnwhiH/6xQauBtMzPRv+vT0eU1iyPzxZ5EQyLlCQbp+O8LJXg/+XL
pxukkg7j4k3wfoSi8zO/Oblpe7+fk92q0WCijIFtYuLxuTJnZGLugkuGCFNtg6W1UV391C9ykKfQ
z/Qc5WxcTXxzYkWPRzaD35KOInr2MOA0XYfSQ0eW3ZwM6BE1Re8C0jkac60Bt083Ai5TTr7PHYco
0xgnqWuwFMcimuJRGAo641zpg7ZhiqkV6gGfPepU/KApqxZufIWTOZK6bCep6d8eudpnCEWJU8ob
jxhcsY6MDNdh3y9BHLK45a2IiOuvFZttTrzO2+FGdLwgAZcVSknNhs7OskPZxUt40bjWRzkuDiHY
BtxCs3oXn8UuJcU0k94KSY+PbVX9PrFhBt4rYp7mv2X1VclU+ZmLVr0YkLh5IbVYQzs0UB1u6WiD
DgRueK/5FTrGREVP5jBqSFYhzNJ8x9sxamICFuNw8Qv9hR4VGNJc+kPU957TVwAYAz0bFdKNzwXu
pNDdr/k0skdOg76ui0dFS2xOqMtnPlOfaJ3D9yBtFfTPKkEYlcUUQyGIJx/KCEbwJRqcGLB9Kzej
7m+AUzhknUc7G7zq6UDMLrjE4qU13ox/NDCpoeGTKtfCPJ9l4OxI2SJ/tNxQJBWAJgJJw4TbXuwi
aRqqIzqU6EFj088uDN34vP2B2J2siGYoG2NFl22IX9vSGrXZTS+kLspBGr/eAk1Of5PSYaeI4aws
2Lrg97pPCHyoNyGZWqFn7kotbU/u4Vd+nI1ZI5F2OdJs19I6VcJtqFwBdpdypRufa+kalFJs3b8K
7NkPf6n6CRjFqtqQdL2kxDxtDO8ze3SdZuMRS6lpNEt1hBvWTwS5gIgdrus/JCok6O/OfuXEXXlC
YrGefNFrUcPWIaMPH1MfjfCCi6qL2Ek4M6AppI4LjARN/nkEEkjS/vNQlhYJCKX959tbveBu4QV/
QKcmGnyX/WVyDQHQTyCh70XItp1+Q6DC0Xe0Zze45+VUQAMYWumcX0U5LZQhO7z32ZrNpww4So42
qzS8sGOLBumiVVdOFWynmTq4jqz2y9OMXMGAFL6q2Gfnc5j7ab/eAlWW0sqm+HEw+q6igYB94khT
z0nvJCaJB0xS+AoYdlvskR+mXOMCXJrJVFRNJ/V0IUpH7Peqc6hMQx2il30dqSuok+NVUVJSjt+Y
afF4Z1huT90tw3mhGyRHeJmIAEOLtQWDER/1JOJ1k/e3F70BPC+2k7Dg/CgqWs1WJhs9wQub+GGL
4st6oBLttqS3q3aktHLp8j0TyK2F3NJtFku+MwQv4q+/oqrT16TbLFek9h5VeZzrxWuuBGoLGUKe
RzUolxGV+Nf0u7PxvzZ9lcaF0wThukm0CYhXT2alf3BRdy++NnPRnL24D6+ZykXREKg+YR+a3s7V
YSlvTvv1u2XxCWq3LfMauHsGw18Bo2mkHlGhBSiu0PldR6+EoxuWZ/sj4r/ZJ0kF4Znd1jAFz0ze
h8gdmJRHBXOMEdxtTcf0tgqCyahLQG7a7+w7rvA0qubgMNRfAKhtUMXQ1LJCtrWxlXwDBLOrqCBP
rJQzBdZZUMBP8A4zfDrcMQlVoSD61AAeF5f/G1Z5kuoD4mCnXNQ6hAAFiyC/vyDMOLbF+PBHvOpK
+HoRIS/kv0v79Q8QbtVHX1huQUlhUvMLKYWt0KiZrc5bysaVv1Uvklf4Ee8ncpTr4BEvv9RDryLJ
R2n9KOai44sDQHmACNWg7Pc3e+jdXZFg5m5ThfO9FmPPsQBZUMQuEcbZTMQLuHnbIwIJoXAFq5dV
TJhMu3wMw/hq75hfvrbAE4tt6omf4VUQYHhVybEioIyDgKiuTdRgO/YriXZFvRjC3OhuxVYzFmN0
0maLRcm2BKXM2tTuw9elozAH+gYENffMiqHQ5Uia7/z6YegpqKF5A/uMU7RtEkKrWBBma939ukPV
7KR8t0qqrQd0KwXR2Pvxx9VyyOjGyia2CLKcx4sNoE2kL5vLxyjRwnb53G8/UQ4lMxqMHqw0uK5V
tD35JNyeKScO0E3nudn05Kmg8BCedW4V0GtCFf1WO5oFvSHqcnTYTPrrBBsVvzZIhpbt4E3ZULLs
2lf/CRQ2fnfXWA367pukAB/AQ7A+L2kdBmOWiiELa1VfiQqzCfmU1EV5C20al3IEmXAYVcDGZNu3
z4m66TZvDiO5I6yaKyuVwfBBz9s4L4wxnWlS4tEY4D6JwTICMqSDD/HWJDxLaEXusuW8cCW0lKAM
WSyhyPu22HunKF02VpO4IFcAis0I2f2G2iQbeKE2j/JZUgonv28ezTyuUV208/IOQo6SwM3XnRRF
Yz2aO4Imc+BKFs3cSS6pqYCnxAjNqHjUQyMWrmd0WJu0wkoyf8UThGWGOh/NRgdNukmz2VzHsDvJ
w0LRrRg/mdBRHF2+IkMQT4Rr2SaSAZJK2G0pi7fRlq/3gNPJFobUyAElhKgY+7WJGPLS5wDOirbq
w3r82e5vDrjZfuxj2BKSfkceOQHdY03BOoejFUceVp8UyLKAYJ5iWOfecPT2qVbdErg2kUh7SUH4
b/DC3+OHJg6pZm5vGejH3y4kP6H1wnnifG+NllHBH9TgnvhRuLPa8ec/PO25OOBt5VaqK9ESd2dn
KycTuUr8KcyQus0DsEbWi16byyCSQgl4ofMPS9m9+eO+qHu/ind5EAh+vL+vdjVazfGq7xg1QdhK
EzA/TkdjWjRLcmbZ/CWeOfkoFv2FJKD0EG/i/XabuLC8leDASJg2xEgHjxtQMefNEu0jg4R6hmeq
tmgXelI9zVbjI73w0C5uk2/pu1cPIJcj7Q6jlL8VZftNxiAV3Uw6I4bFEFZxMfz11i1cJJikUgFK
yaFVaCu7xRDBI/DM9jSzYfM7IPmNzjXOzMjsVvIZUs1DnyGHDpL5z323KRe40mJndxMewZsSBO52
57aG/ILVMiG4kDiJpMuRqz6N153DW8cT9TgYcuwQp+Qr/AXQfy6UXeAEBRVfJ3eTbYOilTnt8izQ
73SdhIw+H1CVs8csaoC5EWMsRvvqE9/adlcAW6bSeKqIXD/vXFuJY8Drqb096aJ76ReiyuOsVJCe
vd77j7tJ11zaA22uhBTolnCO8JbiVwGpfTGml2avatxEExPgfrYvKb6xSLcKJwejIVelahWfbJEZ
FFP+S0wFCp0LysiDcfOIwEStTAiUIUYYWa9M3K565WidwCVCLNVTAXD6cl4Iopaxy0fhKCixRUqj
LZMZ6cIDpGyPR1M8K35FcSBXCU++HDtpc8K529+MeaiWASzJTNzYgGsUry4NHyD+aTUqOCdjKGSG
vJ4t7Pu1urNhILvp/sNF0dPGE6bGjWmsJKWrSYBebW+fddfJjfxMsJsQBL68axocqdDtQkTDXbuz
uHJqCzdCZB0i3zOvPs20P2jjVYYjsfxDPn5ACFdRL4VVTvpoUNvh+0AjRr1dijKEaCkZPCLuj3Hi
mePPOR3HdoMVzUh9eosHPDt0rqTFM4JH0qtzcKfYtuEc/EluEVw5ktpv5x8BU/1XDfqF4pcVoCCW
2y0MXrKWhuXM5cEOPOU/cg1dvVEv3vAXlOr27EukKHhNbm9vKvgqaLSTYvWDZNJUdZLS29UrVrXh
fJBtvZyS0eK87wCK1OPHQQ4/Kpuc6/3EFbR5sfqpyXITjh+npW6kihMgn/f7pRKvshbe3kTXtCOk
8yL1TNxisXS8HY8aFbM10leII4P7EWSohfQsuZc3XC/wR4LIOx5o79U1hLkVsCmkgVBp4CY++D70
W5/zRxqLzzXiHQFPzGTRWHzVQ+H/awVnJ3yau/IbWvbqkhIhf71s6LC6lKWswjiQ+nqkk4B9uhu4
qnClJ9l0sr6uoh4/EDv3zpoOs6r5FgbUsyvjZg0MMJJNd+/KmBk/xPN3Bb4hgA4Ljq5sN4ZFYnm4
lghaZPNkBqtpGLMuw6oYJrzFXc2DxKHmH4Jo0Rpnknq3E/Uy9eAly/ZjCzK6ain/dnlUIqo0yWkC
xZQqMwajilQTY4Lv2LsHBEDtn3Hj6rbJPsNsQTlBLq9YwD/DzIFHVXkz/9akjKpQjKIMCHtVWqfb
PEqSjflP1K9wflwj8Dy4cVebcPCqTFDO8W99yg6cox6pYjEfugHzEAcJjXuFJyXffh3hUyJbIuKH
e/Jn04z8HXCFN5GZuMJH3AvpnXB2u9QLwYvjQbsMWmIgIeCwfFbvMmoA8XRtWQsQ/9eLZFpJRAZN
pK9S1Y1F4caOUH5zCBKuIKmWFwu2ftghxDEzCOZwn9PHS9iWiP0v1PDwKZewuDbbnn03+beCnphT
J0NfkABZGjlYcfAZ3eA1Z9o7LGUTADJ/IqDSbp9c3UqGaBlGrWWjXQrtvl+VnyGxpFPY5lVyp4M6
/5Eo4aPjOWibEr6xAAsS8p4pqlTip+3ed2NiIZ7/RLNC2mEpdNFrgAvHdODyGOz8ZghSwPyxwP75
51NvUvIcLayirSw19vJHVR27XnP9RD6ip91pRrWw8FXDjP2ROdOmY++eCaDl2iXYCmi1IKTIja/u
8CTXiYzF3sId6LHMjTswNDhLhtjeJmzvYMPzPlomGDDSWtUU35txBqH3xnupyAgOT79dcHRo6tHy
CSmLK94weR9kfTGN/lf8XlEUikLFq8oAEP9x8LMZw+lmSGxYRjsVfrBq0l7FflC7jlRkVxkVZkRc
RoCd97TUx/6cxSDoo7dGZnvxNdiXcHOtuCN6DBw11ihe62FJ3w1CaXba2WtanXeZUyVjVyAxOT4r
QVOYMSXINZLiRGyuwYac05vPvMCfQdHwCwvMqI7Lnnao/lcIm6vNJ5F2GvE24I5XEGXZHXnaPErU
rNkO0F+cBKSg26YzIfxzaOT3rVTRSo1br1ZKcS91qRSunKXppgXm7rPMbacMzhoYk083IK1Mk/XC
Ss1v+l42y7wcPZg3zcGuGqtmbkE76+hxLX/O3SE+htBC+OU/vBaWmTMrw7j2Lg69lRCW78i0e8Nl
Oo2MTKvXJgSf5RNrcw/rAm9v0wxO2imctwAHjhf75euLI788EXnm7a4PcMJLIDSG+MWhG+EfBF+l
w+JFW3f/F2FF1cJckmMsl/q4wFtC6fdRg5Qj/DdGHUbH52F76w6+QiRRldAmBwLNiO/8XlbHUe+5
rt7MdvwFUKUChZDRT9ylsJI9/aUW3pzTZSV8o/6DUD0nXvlJR3dzsllovWlZNUh+0FNsPw9pv9as
iNXczILyHkfxlOFHwTqoKffjPSiAX52darsZkOtDhcrHfn679RmZBhFHxjWNBHwSA2/LwrxcIb3c
H2fqi/yqsocZ9yjvQ6XPRSyNQ0BDrvCqqllb40yK1ETVoESkknJhivZ4C5NnZZDYQehgez3qIbwB
CjcD+bdRUmyrmT8s2oiHTTLEHpVbaBNEs0d4wBxhoTn7rFRpRKS8eL272QVkDtGqIbVXzqbdYl0p
7oZHH+oi3Nqu1Rx42jSNoEaTAiDSszw1laC9v5IdguIZTalIxrXbulhss92xZ2dmUz3cZ882ppU6
K0pbiIB/VdNReNzB5dcOeZXgjh8kbKL8zzPBRAmTToFDrtgY3mg6lOef/zcdvYp5Id9mQX5b4JpS
d3uG2N7kAscYqUTAa5hQY1xi8RknyiX9bcqL1djG65rlpFLoixuV/WUHtGfxbnT8Moj7+GuvGZ4Y
WrVhzsTLPWb7vurf4GYD8kjw07iWlEl8bPaAtZLVPa9DtBIQ/7U/kyFY1R9JRa5Gqh2KPWqTyice
VcGW9V6Oe8zbnET6BrpNRjbWB94iDmMBH9cTlY6LBHW/vZYI4NiU0oWobkSqa6kyx+Mn8lwMjVc2
KghcCt47E44kRP2CwVGKs5cF0wwiX/jRuN3ncZbxfwe0bVmmBHyXcAZbuPSZId4FC8v23+P95h9m
q9aCSogfVpLlxCHODzf+WS4RlwrCNfr855iMcfjIMoAQnKWMWxp3qqvXQ+J3l28qwqgK1UhJVg2N
ehtudum5Ft75YPEMclH8J/VOdlWvRlhF8Fki0jqRDPP3pHQzSWMrm9VQYbg1Y/9FcCQUiGdLuQHg
IgV041nKj67p2d3Mov1F1hGl1V+LvfzxuCn4V8VMJYcl13nlnLYktitzq1sxOfH8+5x0AaCgJ1KQ
mSrN19VkV+FBjyf0Mm9kymIpVmJhZXVV3xMMumZcqhX4Z2uZhkUcZDMrqk5MYZMWDEFKLoLShrES
n0L0uXfBqZk61hsNM3Cg6oq2uE4jvAWiMWbeeMffMr2pIwnQwN1YakebEhj56J0KC4mMgEJCidyO
A6X6s9L9KVrjdvUvTguGR7ky+SGODn1UnBRrV7uHBHA5BiAOOwMK/muKYkApUfxrYp14Pui04gYE
RPQDFGgUYQgqGvdHr0MlOEg7R6zALDR+pban2qTpQhaJ7h7vp2fUU+dCTG5pgR47UceTuJx4vpil
sb97ZYOPd7D8JsBpd8A0SEarBeh8vmvFrmEGqL5Euy7GgXLsB6WrPR64RdYYJ4A9je6DL+tu2fbu
hnNNs7iHlI7p9PLhl5kFo8OBu8v1nXH+6AYBTTHW9e4PTiFOwRRjPBE4m7edONHRSHpITVc3ATfS
nxrGBY7wNwRxUyT0FEwduiqbKJVeWVCcuA9ASjnyopaTKHa226YFBNPnuMMo+9U5MWVO+C59lVlQ
xpk8oAoDMGcS1ikkwOIZlCEqADeiLxC6IXKMFXzosgi2VrS70s6H7L4MkEyL4OhgyLTnQmdokCBM
4TIjkWYW2+P+Jzhq2DnJlEuNBxRiHa9W5sqkv6GvzY+tP0iAb8RWnD791F1raqhPposcTO4rSdFD
AG73QchX2VT6dfnYQoad6nPmZ3XvK37VxUdYjfn3fU/lGxZnOuWZuBe91n6Y0NMejl/2iM05R6nr
P+gQ4uT/Sm/lWufzqv+TOYl9mxYor5KtjVSjxkAuERneG5+OnNY5v94LC+ez0pzvPb+f+LhGTV2z
EZ1mS+tYtzA1DyyS1wSO+/LaK8EfmosRR3KGQJgTOtruH/SH1g6Raa+cJ/KZvarw/k5V5C0wXEiQ
212EB2TDoSuTmFnKM15AbsKynq16qcTITKIabiq0+kON2LU9uPSUB667x2rEmxTXakKKKfblnlOs
g0pKVbCWgnm2v/1wQcbZSWgo2PQaTHRzwMWoB+SZZANV90bswv5bkTl9Al8/oh8U8U+X2ljHqVwP
tWejI4rNrctjjgUDcLd6hPJAOzQdC4dKj+9Xa3qIKKMqLBqcHuVezccTXSSmUcsTsGf3SAaPG2Lb
SwxFmQCfInhgVwetra6EC6rMHJ2XtErR8SWr4f6sBvniFM3jnE5FQLpzaE5Wf8Sv/DAn7gw9y/oE
3qwHBXfRbdxQsr54dOWrIqjGetw9yqVmWr9Cge6KTsgp0SkCff4Rd17K3EyZpQ3ts0bLVeJQSJ2b
6FOs8yeLuKLMriZML7i/hiJOU1e12e8B+B6/eXjEzVJuyypAby47Se7Sy9RXcDgNTXvdj1Rtx0B7
UBe66V5i4xbQxWveZxh7PVLHpJgwwqbblUX1EE4KwYFaClFsbQaKQAgpigbJKgW3v03jVxXxRtff
ajGj5YIBIPN7P/9901T7bJTY33e6uEPvpoDA0ckU2uDtHOTef2ZC27b+0SnYJGTmjXsbcyOceel1
4TwxoJJXyQDYuV78yaylGSFjL1AkYJbYOBOZ+Icc/DeCwUxXSVpUsZKfoe6BWmcwHwPA8jP6J7MJ
94EuG5A8L01vLiEdrCOsGvLpMtLnJYOd3IRc+TnDXgVF4zWFY9k+nLmZwuOi+EEbeNSaIIZNqKzQ
r9+V+WxrxmAfkgfWfYYquEGd7YWGv1/jqeyeNxt4c1Yu37Ex3NgbchkPHuUnnkONJVY7QK3xu19C
+zUbQhjZocszKZvwSmzRXSx6gKrNVMjC0Wxu7Lyt9zUF4VZ8bCf4wX5A19N2zZ1E6j37xVsrXnzS
YIWTgJXIchFqs2Dc/u/TRcLr2Gn8Rqu2x5dS6EzbRRt6M2fEPOGgR71q2DXsGnRp2PRHeIII8Cot
/8ZlZzq229/td5nWGQLMh16pwoBBANiFghwmReunDlRwr9P2NQWXH/qj8mlnaPMuqL/iblHpfojR
OHxkd/r92sOZNR59OEtE8fHUEEUuRokh9H+JtY0vshfD5O0I4pQcixSwR+FyEXsskxHCuogYRjQr
XD/o1qD1rDxQMX2cw0LYR9ITohgglvHk0O1cZS3PydEAJ+cMX5cxthxyTC3Lt1mumFAnJ5vFxXV5
oudmkX7C3Ddj/nt7IUmBhb1kToP2tVsIhpj1ZsWemwt0gKkSVwCioMC8xU1fBShg1Fr+wsYmSzMj
0Ctfc8olIV/PSUPCJiQYPkTtn0dFSOIF0AFJQqSkXDuoiwZxV25C4YCB+2c1bJn5B5/VAWrJSQYf
6AVn/xJ1IScU4WgTVtw85Ka3K9eSAJq65UpN7YHxZMTskc8BFyeeSQR1BT1uwbngu8vBfw/W7CQY
T6Ohans/Lzb2Vn52TvPo4lFVGEX0egd/ktDFlJNuZ3+5523fBlsWTtskn8x5YypLkbmqwOxIHh5t
6wpzW8jJ6Rag84SuqvKZCo93RpwbRHLoHCuVSn1QCHkIZpa19V171ydvCXzh4by2p+G6t5LnUxAp
N5movOO8rKqTyNb+XtdmaUeNWe9Awd5+Xa04jE2pMuiU3KThwL5v0mlQ0cxBOp78vKjNRsjRTnBu
Gz2/iB/+M7h4eXDF1Rg5e4AWO/xeWsKsjNR5exBveZLpAcgbI6ttUdaKmqwaxKorrtuHj5ksw6kS
0I54HIK/6AccA0gA7nfbsF3RcWUTnwDowePheTDVKTSun+sVyUUGPHjeQRv3Q8s75UYtGJwtKgYq
u3CULY8hKWtz5oo3mFLrx8RGI/Sz5scIzGle7LM/0lkaobdZFP98x8iKf74uakR6K0y6rQDj/uCP
yP27DALno4YvxwVk6Lj4zrUJJ7yBw7HGmrOlrBId7Lzjh+xXx4wgbNHl5uCgL+EtV3fu7yPxfh3h
D+B4VVHY183ghfoXGIBt6QkFB/2wakSkjQEK3ozNrFWztESzZG7T0uFiRn2TbmtADMPl4Fwf5Sr/
NQnmRZb435W9Jy3mXI3my+Z9xgWNukiRmtVQnFDpD9GPMF8wuCU9Eypac/RVeuBqItVIK2XyKsOC
1O1DlETR2sRPHfSm3VqscWVK9Eg5tPEuya7JaK+Fo6PiOLARd3JCB1zp2btVovvxYbunbbVzUj9B
xY/BxtmQKvleIMCGUhecfXSbStxR3NCdsX3qHyDu4k8NtvYUpAA7YVkqNw4sEdVFVuBs8/82e2ml
Ag/DHcqx/j68eSyhqOb8BkMXcpxHxnTtJKKtXkyt+BYCRaydgL1DgsVJy0Tqt81Gij+ZLpowxlMb
+XpV+OfVQijmUbjNrTExzWJQ9HZ95ZZusf7psNem//GqR2r3jyNQkNDqhEfb2KQkYGE2SLA/TW0l
e8O5Yl1TDqBugQhCZE9OjvDLpS1w3s5k1U5kKvnCMM24eihMg1A7VAnVZMeO+a1NtJBGDv+GnvuO
pKK0WebgrSHJ3AwvUJaaa2KkP4ONDFBfysRKdedTboppEUpwKubF9CK7+qWUJSimdoy62tggPik+
zAEY4XqIteOZyV9Wb+04cmwn4RlcpJP0vfRJjd2BAZFQRAj0rQz1Wj8yBVbA2pzy+vWLLf1QQPrs
8Rw1q6gMBKlFdTJswB/7bzupZo59tYf8J9XQ5JUy4bmmWS1c8Baq4oTdZPm1BYs0FWJDM4NSpavG
mKbD/9VwzN7ihcais2E+KG+UqZvsdEAy0xH6uqm354nfhXfH2WwiZp5pHE/DVPFqxU6A4D15w/Go
ltu64ZfrcIIFeFAmwHHCXIFHLButGLjon8yWJ6UIc3S0kYNKabk7HrkzA1bJxTnYQdczDQ2l+9oH
h8QfbXWkTTN77YfjDwf7yHwjpg8NEpJKV81z0gffQNhk6LUtGES8a7a24OLimk5HDpjYSAkZzprO
Nt5/J+wZEVWf82e9wju+1zTXMSWMPPfKaDgHaLU2pQEHj3jxXlW7Q4bFi54jZpSeAiqZnOaqcoDT
m6jKsN+8IAk+SNrs62Y6CAsUEgumvpDLiAgTOPheiJCetuHxRTdQHR9hcwmV8HZG+YY0tYK4Jrjp
RIKhAtW/dEIHzFBimPfJsAt8q5kZfHQt82tOTc2INNtVmIkHYwKjIVQXv5fNtlrqDE4yZ8Ntk/qF
5xCur5yutsIb8sHc7awHZ5g72+avWyoPlGMvfmUi/PpESA1fOoyYUytjvwOy30PSjTDW+CkJ6VWA
gNK+cCLXm0A09cRvMqhrvs/s2M30gn67yAT+gbrBgYSC20G/ck47CoTOc6dbCTlXc3Bb+D9Ii2S1
0I8xvbzzJQ1p8mFDUMO4Jx921TjYqdp4Cr83+SRX9M3hbhnx7BJSvJxDDYILFbW6w+rkhWHx1xTY
Kq36I3uyF1+pAJmu/XxK+Gwxe1yXzZkVmeq0p848hKXRD6d5gBY8AIcFqYEy9YOfaJlK0J/BhTX7
SokCIOaAgVxr9G5cJOMG+6pJfEtW1fQM/8S827Xaxp50dcKOZCgbz+jzJI3hr9/TX5fsFrj16HEH
wVLfKz3F7WBJzRwoBQthCMx8b90b3+m7c6s3DEg4ksExJ8vIpkE54TwneHX9Q0ufFqjAeYZVCW/G
v3QCm25CwJjkRZVuoJUNSl+mFtUr3VITiGJeEsaeyf03mXAK+bo+tfA1a1QgfguV5J5XXaciBgbV
NwdeQ12O1kS5O8mFMwPsuKIY1pX3r5ENt/4aU1+kdDxAOA3xaiUdAsI8ugOV/ELYPLu2Vd26sTFo
Z70WE934b2IODftp4UC5JdIkzAUo/iU9gVizv05qv0szUwso8U8vF0pul22OTm+4XYvH4K1g7Xnl
9AOq8yXcOSBj+I2xUO0G/931T6VdDGpGtCENnnLJZFq4/EJJx922GTLiQvR3Qj6Ohu7ps6Y1LfEi
va5go2ndBjg03XoYcseDoX6OcMzzDfG9CAqG6c0/9CKzNW6691dYUDs/mljU40V+CdWTACOYKoug
BMMaKpO+s+NmBZrX3AXysJB7VnDL989p0XchFt55A9j4ShegEOzoQc5/erYT1hs9yyh+8lGmyHU0
YMmtIt+dBC2EqQcC8E80Yrf5rYJ0iibIt6vVlAmTsfMLowl9bB+Lx5FRZfrCmp6bLfZQqMjNX6dq
+aASNqRzMJvzAzlE8HGgsinQ19/qmO5aqO32Z+hCeOt1B1uptHFlxEkPWR45Ix527JTnbnPY5L9Z
+pz8KiHF2ZAE9ujMVHrr+t0WT2QTPVt7O9+unyNGcqwQSMtugtnvWHtooR1Ay4y5SZbF4hzGf9H7
VPoa8zIot0EhlWwrU8b+PzKwYUQHcFGsIR22gMN1TxhKNOxLMjHhwzgklzuw6yWQABcOTepDmqd6
OjmFKtgsFQ6rog4KrqlzlyhtmuAZuAu5R2+pvTy6a32SHIL3iycva+73J9PVG3F81g1NbjulbeOl
8DIs7CdadJ+iT2yr3P78X27q4UoviuA5eLow2nZVAMRjmf6uxB0zHreusBfejvhVKROZ8LtQxcvK
1N4tCowCYFMdwa96bIr4cJ84lQzsoWTwTXeLcI/AUguJyur+WVE21BFpic0b6bcCrl5LWStNdtpi
qMV2CyU6/q44nT1790J/7+ntiLdMRjJRCvwdXsjS6nWVyEDcXTnPGbyUtIiykqzFpGfEhN/Nux73
f6/UsoNoqKXwEILNlIMcwoPDMxF9EXHusN1TgtlQZtbubRAqZyLDDT4xkoklYD+NpzNxlXbuoY0U
YcWYnxq2oU4Qu1haf3DqQXSMBWKXzYi2m8yGitxmEJD548UAk/oquVl1C43vTbrRbjjZC0pabdoE
Z7x5o0Lxdt7CkWN19nOqusmauHYqhL8+E7lWA2r4vSI2zq23csoT1wwjH4O7ldl3hIJyPSRB8/6P
b69Vz9qDdbOJY38aSneTwq4gft+4Om4Ljd7SZl8p09ccBx8b552mFRaSIYwv9HjrmCI62UQbbL1m
D6Kuhuqi7AaqIVTLY+vMKu9vUWdUMCMCsMKNS4dj7qFL+UW5JAyn19EDnfCzOmJXPDeezaK0IzTh
Vzj4tTdeaEVz9nQmi8dd59V5zku99HpOyh2RDGDtjKL5IsYgkg0kHAIE5y7mCzJjU05z788FvzOw
hbKMCCaYtv58zmXtw5i8nN1MwvoIJ1B84gVqZVdkpccLnaheHXFjHtrVen7tvpUfMC6s9XtHFuFT
6ICR7bDebEJzUxZEZqMOyE/eXHp7P/YtKVg+xwBnAqoD+O5Y+XJfG/aIVDo1JKwCWs4dlFfOXcMJ
sQwDhN/yB7oq7MabBMHjnrbzVfA3AYsW/iEyCYr+ODxOwjibSSS+vT4/uJx2wFtKT4+A1lqy0FIk
BJvP2vHa/uSVb4OdARWc2/eI1Nojf8iEz4IDz8CDb1mMnM6U4PgIADLsbCCLNjRridiiKSif9NCp
dnM+J/YEN+tqZ+WwwSlW1ZBxST68upeBzyAPdqd8ktppM7zf831ob5tPgtNuZ2YxbcjHV6uyPV+h
G9bxAOgxD0L8RmUPWP3QOYTclcm83DIUCTIi7Sl9grx3sLzCAWQTKkhmoHMncYSfBL/vm8MUUbcz
a1IHbcMQMdo5NDsfxJ7I6eh3U9gloGTdHVnT5U5zJtfSK/z7dku2fLjAr9jsQJJoLeuJIBx6MOXy
cMR8OQbGoCioPK9kU5Xwi1YaLcuozuWbUE/7s/xJluzcx1jRjkbmq5SloFl0LF3B17+aEO+iF1BN
tg7mswbHrdFoJLzAX4ykhWjDW+DDpDlC7ydMDTC6XdMpSGFihluUcrjGpwCspMx3wHmG0fGrdtY2
OmmiEV8kNQPsr8g+hIjEwZXQx7oQ8tpeTW61VE6jRxUZQL8pvN1k8aLjbnKrZ4kS9cKx2VTLWsLJ
a46I6oZ2UGWek/DsKK0yLw2Gzoa4gTIUBKWlYV35RRDgKMB6ZUn0eDhJFZBRmZ7pFA/slWvIqkWW
WKy70mHeb1+iUyrg27cJ+LfIs8Nm7toKWuiQjsc6jGXKHZkG6HG3bTBehsdbkm1uqoo25bBOooF3
bLwuIg+9Cv27r+lyTAhnDOs6DcKt6jDoco1mRyqyQzrnPy2pOi88TUpw9eXu08U/J9p/jqDIL8Eq
csVRD29zGpvcnGjcM8d6VCBXfzTsrkT98+eVSiWNi5tVL42rX6rNMd7nvN2/Qkn5xw4GyjhOjdvb
vgTdB5gZpfyUQqwyGp8+kPvFKcRT5RecFS/gs6gnTJ/8z1VN+Z5X1aMkLsyBFrXEX7WpcmXJyB49
Qyz7jvd/8FTXEPmpcA0CHhJIpu5fLKG+hx1F5gtxyJXbdsSRfMXczCyO8Yr8d4PL8iMtcZJisyGy
NUWTNERBGF8oiMDlvHGKcpMejXDIfOxD7iMgd6a2yUvJUB0sJYg4q+2/vTA0lt0+g8aDtEv+02vl
3gNTwDogZ1LlvboSwITOVf9Px7Pt23hwUUveSRQR/wB7b2Vruo4ND57pYvY5yHHReD0FgWxbHig9
ttUgTSB7UYALHweAoMnUE8m3OHxaZ09SqPLXmRIDeWPmbpWXzbiZFWEdEKQwPNgLCvZuxIRg/BNd
vlLsQ7IElI/y6jba8RCGBS87nqVrj6XRH4GWnSoGnFSSwCKMYIjQhG9bW5rqji9PtruZGJTzX/eA
ewmmh5QFKfmVhMlHRaCA4+FlF604JWUbmBVpF3diGmziUHs3YsMfexbuiUV3dbU6/XaKiJlCLFRk
PhykbuSO2wAeC6ZYjXEPg5GkDWkZ+IqQx8rsRk+itI+Lo7cL0/M/ST7GXcv10uzeEdl2dKxfcruM
3ggMooPdadxsAHzBhueHNsE+yuMTPT4csoHyyI58yu7tEhoEO5ph5W/bjmHvmTH+79ncaZeYXJuJ
YIFtHnLc6Ykk2mLWonG6vNF8DvsRb0XSyM/uwrWkzQKM9jxPWU6Eae4iChtvL3TgZ1Hpu3yQ0kbi
llyocM1XQgcqY/BQCjc9p+yhO4n38vGzVlZrZiPR3kXrVZVaib+5d0+Nggq68fxaYnm8pceGph4/
okMWWxoKEbQ/lOyRm7z/etnE+fpVdGh8/CMc47CSyqqAS9g6RvG3EX4BMNY0Iczi09aF0cN62PK0
M4ZXSurRDu4NeF8cBtYlF1k/aajDYDRHkBhfXsqM0KZVPj/WgjLmI+K2SWgS6rfgoQ+Q+wIYFXs7
d46ckr9HAIbBqgO5BSNNe/xUkxsSpRAYYNYUgC+zvt9jlh6MbE54pLjXcYLnZCTLXRzFcIUNC1Dh
uEkxZw4ALCRL5JY9/u+aLyzhHgglIpDttTLoaQpBn6K6y6SGS+f1aGCLDaBM5zofz0WlmqbMmiST
W2HYdvxe/3xll7yT4Ecv1tZLwneMXcPegtBGqc7xNND3iCVip0OXl1U7JWm8z5euLuIycehSke0l
rFfKDFqwrA9V9dNYUAdTR5T+XpzIP8ntI1SwNNTYjtbVgagt7G74Fx2Eq0KmN35jxuFOFVvq67wJ
g8fh4lm1aVeWGpW9FPSzsxcN1x/gD9IcTiTDXkqiXjaanTHldhZ1wXFUxq7aQu8oWfd4kfy11WRu
ovzFKgeahhv0Qd0eRH5WXEX0RUemu5PsGIClEbCvSkVCxMq69naEVIV88SJHjGrzjDRVdrGjjMmJ
CC16smhzL076qXZxe1yMRBvZmkiEniEeP9JwuQjP+qKTH0atLR2pP2rRrQc9YZBc88kgLZn/rCDP
ie0kapzvKoFXNt05olp5BqZ9XsXwOvhfhzQFk+evVDLVgeSd+/qhtj0tIexnLVm5u3hAW+B5Tq0E
CqzZKTazBzF7yWOQ5bYUNY+dhxG4bMOo+xvL+/pdEo4fEvHWw8xH6vXRCaUMDo/UG8sUJNtCbc+h
Xpxxp6Y7CAGBdq7mXiqzbaJ7wtbvJN04PFzkOiddyILN8NconjBxpl6KrCU9N0DLzLujIW10MIXx
BAJMGbLL5YJBo8c3lyr+/EdGOn3A1TEGaHxsPNhbdC1x/utfoBGVsdwENfQxeqrXmL/1cuoCgJTk
VworS/TLX0YsLqkUwkLQ8sRiH0HHAPlsPqq+pN+QX9Aj5NRTPe25OOs8cIGAFbWs5FnMWU2wBJ6H
qhNAl127k8ape9/OAtFxKfADRAZWabNA/WlCTZDGzjSoQGFWCD/Ggmg0TqecTyvgz6Cg9cfQxNe7
DaMHGPz1904KhVOypRCgVUpiEQAYNcXf3A3D9xyUer2dqmIn1tMpMAXILNjABvoroht8mNfQLyio
sNtT354s2ZAUIMPPtTvnZQswFwGdP75jkDCvD2eULCqLJXSevpXMJRIszmBEtBTBEvw22W9WNDfh
4ZS1r11g6cAQ8Tn8BdoBqE2QdxwdgxktUCedvSDC/qO/PnEYLLnaeVLSidut32bqwDi8CtrcoCpX
faqcO7omVI6SNjkyQ6XQmGfW3H396lBfbb+E8JiXsLdh/hq7mC6cA2bGd7uEazwS4nI9aTL917rs
Gmssln2CEGlvTcyU8WwgZXbyAC2bHCvWrXTNrlIH2/3YcG0a7gW2Y45EDGFwMhhnKX/A779tkTMz
PDiZS6rQ0HBJi6Z5q7N4ctUo3y2Hj7OJMz1perHFNcfXxKp0jFQMvcMvfskG/yBVsxw1Aq0bBMan
kO65T//Q9j8pLkV9cY3vjOgT9IiQmTyMhsZmlnLdOs7qZu5AzkBMKosJ0Juvig08e713BlhDIb7K
pMUVqB8XAp0JvsDDum1S/fGVUyZ2OQJnv3dVG3hBZuylKbEyWremxJZEUuW5Ot83xeavcjTlb7/s
rz/V5I76wPxnse1RWURBK3Oq9Ai2fO/OP2Ds3xCpr4GtWTsdmhkeJBGuhgS7lFG6w+kUaqj3V3n2
HOrP8CsZbQ4Ya1M9m2RlLGOVRCNMXFTCPA9iEFnQ+k7h9BeB+XmbqF8qwxgrKbZN5BURL+v+qMaH
dkF5jPEBgrWKCVmqt9YS9SgLz2U7B3ZTRs+Ap9UJedbRalzRXwEaatdxog9ED91mTuQTAAVNG9tj
xnovdbbo3Do3yDi4MYW6lm1AXYXy7aJq8oZ+wQco3N5bONokgrtQlKCVjuU6cLgoV5WX4QdikBOv
AZPuPgChygkgtlFCCfZIpyXrhBq9/itYRf8AQn1aKDGGzQpe0jS4S0jJPGofd/QwT0UHEUsXttdV
BzYxe3TIxiLs+eFhRpU9m7WRdfRXUwrpYyqFkipp7CvNvOK34x+sxDLG/OrgE2q7UUAnI2AIXa0T
aUo0oMMzcCTv/pkZH/Lp+oCSDDmxIczEVuqFV5DHGi6CLfXbliTm6w1Hq3X9lPVNfhof0LU1RBbq
Zo9elACrRHZysA1auLikCJzLaMdaTCez3q0yHmMMSqoHxDIZ0QE5A2QASRC6Bi6lDChR2TFpKSGO
ij433gnayzqto0UdlEDckE5Z+iQvxO6OhVYnkcEKK8zoyO4qDfpn/LL497ZrKH9kjW5u8d02KJpL
oKTOsMI4RQ0OSOCldZisaoUZ/APEMVyDyHwBEznSXgiJq8aVjQioXWcPZ+lOQH1skC9TjEy6uGJh
JJrtlBJQrYjcgW8kMDDupXfBFcnKJebl3WODtb59k8MFmmG3LZK/8XmsH+0HlYpKyauL+yPSfEZw
plDGpzUucl7nS+WnwVc6RcKgy9BsUgyLiN3XXun1zScf6Mef0S7xOO9JED9BfqUxZbJBO8T+MVEg
ox9F8zJOmyB5OikSSTjUvQTJUadq9JaWljh4XmwemTHUs501E6xfT1NNqmY8O6nw1xoxKh9V5irJ
EofCh65P3kSbFq5D8nymUYMPmCqdX7UlRhyD3EpoOyhNjvLvj5EeTMoj2rBYDCMgWCGk8i2ROuoK
i2xVtpLAVqOf1XnxEZxfmgfU/47nVvrYb3R0CPISIDbI1yW5qCeR9qpCM5RJFbIaKS6XnboNzFNy
XIjuKQ2WoK+dzmKCgU3vJk/f3WNs/W4Q7gHKY0kPZRCPqn2VjObtKQf46xxcDspX8hOfVyoXzwvF
HaO1jVoaCWzpfQZ3RIdxVCnAgBuzINgjzvEFJ4Aore8kxGa0Ur6yNApp3D7rb9WRN212iLhTgiaO
nFBgBVzv3Pxb8EzdwV7JrZJUi77VpCA7gf53iXfrdedhOZbGlut/hXfMJphnS36lmXaR0qHjQ+5M
y60k59TOBy5hfApzuQIDk+C26XAu50ANx6I/klOAYX/VmFt9uq1KMaado1an9y0dM+YKlC1sRR09
nhMWtfqHq7ThSo/wKM5EsP0gS3ouroocs26ju3PpDyR7J/iE2d91Jhk6UZ0tiHmoMqPatObPFF0j
aZJNfBYaBtpVZaTBnuD9hUUHIaEMXbTI5S/++Ux9rmFNElUqP1KTJeE6uNu9jWhlHakRpc1gooHs
/xq7TWH21i4Akvb7S+UBrbP/x4zYbCh4KTEBx+VqMGhp1nD01diyNrxF8Oed12TqqHtCGDXhh6XS
PpsDcD9Q/zIdxZuIK+2m3Ag8ulvy0VqFIpEzqZO/Rig1T6APN/O1PSP1+Q5x1X0e0vyTkpezu5lR
CScDRLBC6PW9RHQbG5IALcV3Io1I+8d7PoWvSvCCUdZ/qXY9EZ88nxJxLRvbv029mbdB0BJgaA+p
CnTbCqaCjg2SB1/NOPG+prmbOy5L7UjVUYCExsXZcIZ9nDD/4dKYZ68oTrAjb6zILaCQ2PXwnIJS
PTklDBmMYBsUJQ7zGFrXh9q+W2WUhFTXk/8gTwe9cpBHnQ8ok1B+ABFhT54uean2DamGi6Gs/F5s
pmzoS0ChMA5FeGei+QLly2S2f0DHX9phXsy/ep/lrhpdju1eP2+K0aHTIDIMXf+TDLz92xYlEIZP
3xQrmDlMUea96uBC0PUyg3pYOaBcjVnSFPa5BDQCbcA1vYqz5yIKodvwQ4+ko0qSh6lhEdm9qxnZ
4DGjHPJ3hcQocB535qnHQc384iTzaQDQkPZqiuNcd99VqdsZYLwJqs3RhkHOJ5C/gSWvWs63KHC/
qggoNctaSaRcZph9LLgyRC2Cfb55686uJiuajymgvzdtj/V9tj86gSDnwsNy7vwYWEOw6WNrn6U2
VqqLQoURN9WXn2+gLpU0nR+LgHfSmTLgDToEZR4JHf3q/wxm/FZVzKO6Icuwnjf4onQ2HowAYTIB
r/0nR2RSxCcj7xyvKqNf3BuBrnjzCkQobm0SMU/d2aJtFZNMy+GIjPEAKCfi2pGTd0Xuqiwt4KxD
VjByve5TQPB+T3+WJtUUZqQaRTlXafLJuaP3rX9aKJ+DNdkBnm0dDmMegO1sl6KFPKZpcG1MJRxR
RCC3IsOUxE/17SjirkRsRluhyKOIgDxzQAj7DY473025KWKbPmFhYGeVEbGAFRsUg94gdt1/P0v2
pCC1mtrjl9WZejxGPYS1bQrCs4f8G4HWbDvvwLi5Fq5IUXvHNq81w6mvZmLv9ARZPou7QkiRvxuV
EeM/EAIjTgY19wQPjNcfVzFcYMyaB2nQthxy7EMViPUkNSrCYAq88zyukHcxPENoDTkWLHwigNbB
Egl+8mE8DKkVnMElXFbHl9ZwgXZgVTSgzB1wSpfVlt/yywYDvLG8kqqvYz15lxgfu2neqL5qGf30
GIGzcOATv6x3fhTEYKlTuuXGvMD4Po2aDMQM5lpADgTHR5OYgUJUoSNA+nSMzbNRyMOT9sVUUQhN
fOmluj0HhwXDP1WUhq9q+7uZVZhTA4oTjbgsrLEg4ZUYAQ5NqRjtYtdiV5Heg99e1Or00/E6kjx7
mpY/+gvex77zFVe2+H3qTpSj+tEyBXgcdRFWo1tuy1qW5L/LtF9pxbdi5+qvp93bKZ7+eAInYjBd
sIaP10wd0HD/E3zFPhKwWB8Inr6mIBFHGsNLWJl1/dm2J2HtaR8+FTb1JjM2jx9D5LbORpmOEnG7
vV29QZfN/nXyS71Km+1Of2h5dF7/RFMTCyHUekLgbOTg4wmUsNv4wSwFJqynzqwMXNVlS+YDYpeY
f26+7/VKYhcMQZrxNIZUbRduCNC039JscPKv0Y+tFZ05hqC4sXZGRa6Hd3PE3804fG9APMWAgOXS
Ag1xvaDwYkXoUwfP1DRV1jPkP24ctfBUSTmEf9XyOIXbNG3u/hdc/m9qhYe3mE7An4fICU9uMJ1Z
O0+UDvTXRo/mP3ZE7AeidbQK2mhT2XT0sCJc21npzAcyCsa+uG43j1R0yKtOioP2bBt9ZrzsiO+B
Tdj7zoxkFBx1htIKowrvxHrfnAkCHQsrRewcKI5JUfKlkjKRmsfmIPHI2sbz4ZTklOSDAPOxwmXx
VCP9jFIgjce5b6JUjcI1V9DM1rNIMH2hzBMQsbmBXmfMu+dwvguOov7FlwqW1OSuSjTY7jaqtOeF
tmAOO5UX7h2YOmoXDZDOA7zb5/o/Zko5JEOmF/hGhpBcipC+mG4a7f1PjXxXT4Ra6NbuMiQTcoMT
RbjTiE78aTOn7g87UjngN2lmjg+fm9xzQNs6rQQ3fBgbKNWm+/t9HZROjb3WFIP931TSu0f3NWj3
SeppQgD+OyvEsDFfsW1e1IMs+6x7tnKc0MW2Qb6sY6ciw4oHllPvxodHCjEao49THqsxlnfoAqhm
7jRqyW5+jR1LMgIl1mrtyh85Q8lKLSPWfvKwHJuDRrvynDm1j2q9whHiW8Npvg0CzQHQj2ftpkzG
YaW5ZdyTHmSWP8c28e+5f4bHnVqeQN80aWeF/zhtBjqnlYcwJA1c47OXzNGMzQw8vhDqx5pnIb+w
j5Du1nqV8Vf09sxOCOGRZujdZMfFi4QJzBDaBcCI7KfrKCcMl3Lym935QPvu7iw0kGs8rpFF3oW/
+Uj3I/oVmhQxDiZOfdHDK+pLu3WI4uCxu0QB90Rdo4ekV1r7IHCU28PRjfGVfX3ZvJ+MwN0p+cnl
h9A2ZlnFWOApZLqCWTVrxTpk92g4JssY/pnd/XWhNdQUOxERuBf50oURI8HC7dWtkevo7sMIFgrQ
G3AwROyZqeKrdjY52eFKN/gJMwUO6MNd5vjqBbfA7YokfAJ+c7ppwg3W6efygP9ZtLPY+1uCWjSO
hYcZlejM26VZaAdn6AjLRp7HmxfHA0TSTib2yk7g+Ta5xlyoB0iPNUkgIKzk82kL6sE8fsdiuWLc
PohEcNIlKEFho0Q2cYez8NzMqElIsxRbDBNeBv5JCsOOf1A04LQilgM84FOPSZJDy2GnQR8LWzSn
PoYquoHOWiKKKq26fG1fwjC7PxgMfZNZigohIAjnnENKptjLIweH6LvKEAylDYDqPx/Urxw+VYyF
OjllPsmmzWqiVmE9PmiHrhRLlZv0clf1uCTsUJkotdwKkQlUqwleimVm+Pb++LA0PZDQ7S2tDo/l
5RCvK7om9GxB2aIpaNVgVJa6AtmdrpO5jkBCfrvjvNnd4ZljAmFMLrFRkWv3r5+L0d5fYmmz5ZLv
s0vSc7dZUqLrvmwSIDceQlR+jVG8/KfxkCYA+zMj6IhPTM2Ql69qyyL2p+mPW1ay1bW/WpMKYBrI
YrfY96NcH4LSf1/xRPXlCiO4hWOJxmx8AnQC9aegle3/pU209UwtJSi0yICd8FOqFdV/OiTN/zpb
rwhP27ZNGUaFH0uTORp16IKJe5+TJU3/mSao9p3WzNxzd571NAA013U60np+l1tbglPMgnqJZZKm
jS3XhpqjtpViHjj6VJsxDsgQ8jfbdMiAWL9CoOck9ZlsbNmrYucnydFL8HJnmdayVSga6Z0Icxhk
QRdjrdHkvJzBxmvVHGbfUgtInlB7Jj5Db6RNn5bCnpdF7ON9rhOfir/OeUJa3yayBfWb3i+5io7h
boDKEYunur1xg1ZoL+rYuYJwWX6lLQntjLnF6pn/aUYSt09S2B2kY0M4xPz+77D+EvqNSKy73hoG
dqvwrDurs9C6s3XSUBnz0goORXKG/wPVECEtKqns31NcfG6vdsinje+bxXrneibff5OPtT6/Ar6w
6RBbxoYmWfSnmt+6B4V7ZQvF3YSWwnfxk+vhOhLdtQT5vpwYNmkP6wD/LJSjSmvlVJxtLtHjGNBC
M8ieJbSZJv4NiiuskTc3adBKMuR2eXlYTfTbReu16Jb54leCI92/lPXaK+VLmALqnIwy3YeVDHsW
x7EQjcR1vrAanbz6ij3qAsZs3Yu2OOBX+4m9orjzmwCbuNSbtuPxDiQrDKTNGeF5/4vGMU8dg9td
aGN0mLTFU4+OUU36praeyK9i677BYp8RdVqWE8idWYSDYfULJMwS361Tce8Drd+yOpjD+5abxgjL
iruE2xguoiek7sgmNHA209SvfKATCFpe2fMBSIhh0RjjuNXUnAGIITgodSy26u+fR2gLqoe5waZ4
SwBrFFYgLCX7XUdqKWX+4WjrS0fdzOJeAdYkzsuEuySCTHvu17hkjuJColXYn2ca1T4AU+AmJ741
hiUNMEspb1NrKdEUXTjmMFk6NcKb2yQPp66dUh90y1+TOwGte7MUfjA+6uCe1uZhIV+iW7lUcX97
a15jqabTk5PFfVG5raQUT7ZSVwE1mjXpHaFjaluhjs91QmLSAqYKOPfCOL4ZRU/pp1EyOYSO2FoU
fgSAHsokr1f6i1H7eTM8N7quYe9SrkRBaXC2FwdOdsofGJXP3kqYnydSZ9OBkcCNVPdXy5KhTsKJ
Psnge097zv6stIBSiEaM5PohT3DZ0H3BAZXVGyKLaikFXCQ3npSByMxxL6FIpeGjwow0dNl8+/1e
hNjgEZwgFCGqhUQNSNppg2KuHeOw2NKwhhDqam6q3KS9b2pi9QqUeXV+wnB6dl0u5PY+6Tsz+Gf9
kiXwznUs2EJEGKcYS4gXKM+Djky8xVha77qE+KlaqzJGBtVcKUZ0s04uZHd+WtTv+2H8ZRt4lB5N
9Zjhl0KanYvSppZZPb/YpZ6K7bR9ZWMub0V0zm5/REBNbtmXuSM71SXZOatpFwZlnL5r8SSS8eaE
hDzz0fBbTu8Vu740yFlmHdoSgdnq/K2Sr+Qv/r2LE8nhPsrKnKidOrJ8nA2MbKcK7UZor3yBo7bW
fMIB7bR4qV3xZ4UkMA+GFMSLR2+iNNKlVOLwGLDNbjonkgc1u1efCw/AdSfzBg2q+nBJ/DvVnIOw
8Xsg7IW5Hq/ppqK/N/HSvCnmGo2P9rx1Gj0XFNvltNNf22iPlgaX00rH2Lnrcf3gAl8XFQH6///E
KUcIm/v7ZwaVjREuPqPCKrseFsqJf8fvBEe4XD4/IfLZRdzx7leJUaz1iDoDe3pGeB3/gGPj5QtR
mX+te3zmbatyKJ4hcg1ymDI5MaceZVAy+3nQVAfu8qPrqGxwEQHOhcKtkKUaEndxEg16QlzsVZ3Z
RXVgaCGxUcKN0vsLmljYNEGrVBmgaIAIr3nFp416MhMseN18lbkjDSx8vFCwyE0QK2r9KJmNq6dR
D0q8SZJQFwwswypz+GE0WtS0RNpcUcmjJuRg0BBEkHy6UWlfDjyW6y7CqI8isP5nAMYCW3u8Fd6q
45/qWM9OTAHjSYK2CZhxrRuxZfoRdOpSlQ+KZgYC9XXb8eLaULM3drhV5F2/wrjOBe43zc0Pxd/k
oBG+luIMbayEqYg5FlDjE5ITZompBconS5SzOM5c/XAYrsFmbcSpzJX0wyL257Hg88J7BWJ2DkP2
w1NxpMXrh+fN7K/AIfsQRp0kqSjWCr6I05BMZZBWlu0B2CxbMNhgTXU+kYdoKVCc2pBli1qz4ai/
xegQeahg0TtzmvRgAqOnrGs/RAQHuCjZwgZh11UhgTQ6DP0F+iZK+DuJlYtOUT7lO8zKE0QxEcCH
Ylqbzy5ijWVaDSy/VvWQkvQK6IhRQnmJrW1JvoLabVNM9J0vvAiJBzVuESzRbYUdAgk06iSo+WgQ
Ll4adocFHXZ5JcXU1c8mWQIoQl9vZanXgkKgdWxmy6IMpc8dM0Y45ONhwfclKMpr9o8JE3HCvDE+
Cjhspw3ispFdms8Reimy5n/fxVESRDXpp042yWIHrZw2zS7wIv4mf5V6y5g5PPjrvhuGtUKT8Gqf
RJXrfpmKMttG7Mj2mZGJqaJ7NYs9TNrjgm/TV7fT6gU3pSAF/wTF6JOYB35VAhwoCX/9JSMzuREH
1liW1xJ7c7BlB0YPKJszXISQzMUQRoPluqhcpRoKryicUjlm9vrxyzrXm15rSaANJiHVnB2H6v95
catr4zd24ueffSgeHRqzK58jBIxLy+g+B0I81WAt2uLl2ZuBRUl8uCzaglfwypw3Qi0V+Z3vUTCe
ksaI3ziHexfdC9Fcjjn2qX9fcjx3Emqg9x7TTovz706SD6ABw7F4QeA6D7xHsIj2KmGD04UazVGr
3nwRqlAwIA4/f/u5S9kXG7/z/tLq2r8q+HF1Omi83/V9v//zbMfalWp5avfK7eLUcVmPhprbHg+O
yrU1UxyBZmNtsLDPNtIsZq8BlvfAPcrhpjmlGeMJYMDgHshTPepNdmRG/E1mRLGVlRWoIl8tYqAh
Cm5roMXHjCgnMHpw5U6gEVCHXChi7gZWDE53AGRV8S1T+bZU92cWX89uEHqMDHy1mDJd+3wUTo+4
plP23b53rVvsojj6Ckm5EM+BHt44F4gXvtFWX8OoMqPY1gdK2QgTtW77XPTUIgMlLI2ly9PH0Q/r
8hkW44XoKqy2oGYZtSHTbKViq0zI7ETXR2SJyjIRLAA6oKsqrQ+tRDdFLFn4EG2Z2vj/jLyNmUSr
WUqCuEFsLFHA7WNxFLeloo7g/DcOXMT0RGlRnu21d7mM9l2zvmOQlQNJznU5WDwLjgSkdCXBHxvb
NkiZt25KRlRTQpfBiUB0uGDcGpjYuHKxrRQFPlKBzL8qtGpuRVUSoLpM4RKDN+NMLB5W4UgxDPFA
BvX4nfjnwxZ21tpbLD4KjLgIc2Ok+zvGSv6olvHNYDjFin2HxWIeXEOxZouweDb/+L53tERRnv0K
0PgBBVPJck3OEaceDvlxjN4jejHfBnokZDLxsmT2rnTUNr9kvXKobfhOC2sbpKHYfnpF/Gep6jKm
l3gx4NBaRExINisquaErwoXKbZ5sqnDSToAThu9JDWoOIvSgfc8ehrxDjZfTr4QqNKKqXsn30H/K
AdQdYBNaD/ciPluGBKsJG9NpM8bOi4EPQkvPvvSSzkNz5sGJaD+Exw6zJeq66nxtjiKIHbrWRod9
m5Y0L5L95jl0gLrng2IOzbUj8pYLkdNcY8WHwvg0s6CYXMajaaWlOUo5WU8mC6sk570cwpxC71Sq
yc0T1mxM1ziO3OJ4U6ZU1JWlLBvXaWNRvS/QzIberVupNSaZ1QtipZLSGskyH3evY3YeMyo5lnNp
hTel69p6xw0Kx48m7wWWno2p9I1YqQRGm/L5CuMKUMclfNubPEmZAeeNCKGOKcviDtxziIklP8VD
Y/Gy0/tVQN9I0RF+YkKjFZGgmzDGg/imFZHTND+wG5cR+Cy4jRZUnV6yQk4vWtzJnwTnclLMf7lm
ddbtIgKwB1ifV8cO+R4zbIQ8au6BS+GaCrppxNMmB0oScdyZdk98NHx1BCisKwDlooaAuCrFqhd0
6N3mjCmkcIEIU6SHV5tAyBjXhAXg4nD4idmGEnv14hlrh+P1eJjP8GNox8aoqaS0VKprperdquUV
hobylwuE/F6npmpO2oulD1ysCQO8HSCPUmUxjfO8DxrjP8Ne2NhG9QbnhPuSJk2Y/TsX/gbVm4bW
9AUKoI7YsWe89JP7EDQakwj2YjFKnZ+Ye+vNY7FcqY7Ew0OwvDXit1xkN3xAaNvlY6pPKzGYFu6V
w7fngXKlnP3/ZMK9Xkqbwm8b71D0N+WVd6ImFTvGdBRsrUuce1xltRJKzeyrjPiMubXo83EZT0lQ
AHyLG/bgk78t86LpkDjI4EqgZ15c6rYYDq86r++8iwMROhYPW8SDy6cE2VhsTtdNZI047+R2yFx8
dkE+nxMNWejerOZiZ0DCu8abK94xZ9YMo5IqOml6mZZ+Lakvb6gVycBTmrpr7pLMBPgTSvh2tXj9
+nW04I5aGxvO95Rx9Q9WmlGZbim/F/s+obCGBweicN7EiJN+Qo6rxSzPsV/pJ5HRuFnwXF57KHFU
AhQ5JTF7bHFUmUamryeTR1qUUfk1RnLLKiizq6WL2+IZmMyS+4cWKFUe1eHP4yyduRjZJqp4ed6z
rXCHmFaOoSq8MobiqNLCyw7Nplxg8jWwuIARL4VdlLf5VpI9Hx46MLdrnWcV6fRn4mY5j1O8cuXQ
PCqLHglr426jPp9X3Ax1VorQ1EhaH1D7bLtLPaYOo60bbSpOvSUlSExsdBQN+JrxHmoRcPQasTA2
BIciubkPqvWaiXe+7iy0OZoGI159+pVFcIr13d55EwaR0UyKgiMgsjX0VxUggzXe5R8YRHXAubAY
YuTr5A3uhS5GBOnFajkPV6y4+l+PBgXp71+dslrld8e56lThKP99Qej0fuo3srsz9dP4xsXjyBT9
SDtmS8xW4DpBNrvzzgqVu4vljLq6fSAZoG7kIpEUgATExqKtl0cD9j+gxI765RLjDNKRJd13OrmW
MSzDeEL3VXmeXX1MNeIfUYVkj/nurf0ab//wlw/ydCHW4L061WOCYovqRWrCqXbTr1Om4zeNHV5U
u0MWdrFnjZPV+CzPJHGL3CZmUJV/j/QSbWYXsIFodwCGxoQblL3nDb2ATgp6Ell3iNSXNwARnFKH
2N9zfrmAIx+Tkx+0oJwXDQI6CyTFqVVMLJW6qnIijh3DsPk6SVISTZrxw0t8zME/3WY8s36Lur2d
Xsk1P35hHCGaOeOC1TvwmVXf5whv/PZoEHj2wxCkLXdvnvXVsGoWFYmMdhb7vtZL08wxPGhNq4/w
5dNHNFeJHnAuMfHs2FJtF88J++bhKUZNJFTHMgxW5ATXM7ePCahRGXmP3gMY7yf6BiweYCUey9N7
K5KOnrDwD1qbcAb07sBUkiAb5uY2IljUnAI+tKqmGbAqImcasQ9ftrZg5zCxoLzSBl3iXELEceIQ
Z96RoBQsg7k4c7mjMUrIa/qecDjQRaBX7YdlqcSvUZmuUE7IXf5PmdNOkD3WjylzL+WZ03zmJkYx
JgrNNxOi1UHqTeuQIdVp9Z5rUe2h64VtjwP2oCFoxeWtPzWRLF5XrLkCooG8A1gVEhKxI7c4zpKa
odNkHNrHFcGRALpcQyy0o5XijaohiiCvm2EH2tyt9/Wxx5Aw6UH6cIqHRFmAOOfhIALpwZ+EuVm9
3G+RxENFu599XfCQKTKPrFSb0CsfBjTOPiCnJpsOKR6uGja5Ui7ayC0BeD1BrWnz4J4CAy6mg1QV
npF0FSdwbpJGtfvhSPrAcGJho3+YxoR1siaP1soYe2Bfvn/JD3e/Zlyd5y+N+CtfwK7lQf0L2oCn
RsNFwQv4WJU8I/EA6CcF+xbGl3sdLwHH/epGGHHhdQkc3NbGz1hWJuBCIeMBe/of9tIZC4LmcNw9
yB6aDR7ppmXHqojdnxAnyPma3rn/lknXv4bvmAE2cIVZr2gxv+tsfrRtrA9UJK1jA/mz/Vw1p6iE
5TdUP1BIKFI5rzfdFvAI57bMuGA2A4rWBYzq8y6JPQfK9d1HIEcopwG8UvSmx+WAEwlk1PLbK6q0
Z56KJZDnUAoVC/nStn6Y0gLZ9itFzfnWoUDtrFLlg2CMZameVXNvCSTRPFNb7B3DzrvMD6GWPBnv
5sUpfzOf1hJwusHOF4bAgDt/y/SrV2RHT2687EUG5va98R3sp1tXb7us2u4aUd3YFwuTQf7E1UJy
5a1Weeu/XE/eWRwYCKMhouyyMNBXhV3xBXw+4oL6tuGcgpTqxj3af2D0YDBIrCTI0q8IGuP9SJlR
SWlg9luEOtYVcz6+3fJEyvSGU87/9Hfwd6y2aKUD7Be7N+UcpDvnvdBspanNNUa0fGH8OX4LGC5/
D/SMP6dLl+gz6d9p7j3/kJlY0L1qFksXu02B1DavZc8IGXZGQVWntCeXBX0yNovz2M+DWG/uBxFr
3Akwh8cZIN21giVusTLTpXVJyt0gXLCunsUGfP4Nksjce/L+a32fh7+nEyOLQCmlKcFc84iM5dIu
tpbifTKjQbyuN+qZZcV1hJG4A3ApUm1dXxJE20PKh/P2z71U3Z6nFRyko7YRuZNn59LolV8vADm1
tZuDajfUGrv8SNfJ+0hw5mo/rUqe0w2qhTetGXoFQd2jY+I240oVEfIscOD2KPpJ4alXU9vU2iyu
IlCXHtb8hsKsDpi6lgvbkhcJiAdeCeZgfhO2Mk4Zhd9UVYIfrYFnVJIE5lkPivGaALo8VKDUIUet
AtSYrGlg12ncbW6JljzSw3o0AQAVXV1kE4G7Q5I5pdtR+XUMt2JPFRrE15sunxNUGSyoWeNxwie9
X1FdRlUYMR4RDqNpdsbxmERuzEFNcXR+cS+5qXmfUwy3HOUfNEKRHUr89vYYyq00TApmRN4iDghg
VSkue7Y2UUoNZ7UUjaOgKkFsXL1SATo/wpPwSMbuWxYXNcZIfQOjHEhor+OL9zfVsHBr9CndE/wY
uqaTM+HKl+ma+VGwcncUW0oC6Oj/rNk2cIIR2cLvBcOW8Rysy75rFCseOBWuICSAcIqpsahYAcRx
lGjQ4jeunyRPYvFQoncFesfopzpbs02huSMiftWm3vC+uinv2IDP7Dntrjo7bcTILu5WKVX+HJcA
4EZOVb9JzqA9dpbGOLKgqmQOU9M7tkOmF+mUs9080wgu6lZMXenMQQo8HnEzSgd2R468Sz51CoKZ
euE+XuBOFzGCPkgtQbRFuR7+hbMg9UvH0zBW/0KAHbc2CReJqwQNjd5vp1zeYt8aCGVXE0Uq+GAj
XsN5YWOJATb49nJxG/Cuad9UmDzf1sPcet6IFLt5O+f1NsMhaAzdWC6XFLQIQGekYK+ALAmCp1fT
zmSBPPv5oj8IOyx3w3/T0Bk24W38bi/GGjVZdP6XzFAV1D7Xlt79LeKhvM+wcibLlZw/styPAYfb
01skKdO0GEcrTcGrBu/cKmyNdIXGWDKDzTlxy1SwQcKXsEGHgdybph7MEMiAO5Vi26f84wtZEPVv
50Gd3kXC7MG/aOPEjUNrI/CwZ5V+/7xUeQhuAyNlkUH7iWZ7B5/8zTEPFdKao1mNKy/clAK1nyUF
LRJavO6dbwkQO5wX34OPbyHxBFvhpB6l41SSZ15XPL/ASGaM235iaNvhqgZoE08M3nF0nDizv95n
JsvKZ0jcXp5r0rTi6BIQ2HBiwqQ2O62EH67Bp7wqpW7BbLO9SmjPx4BvbjyteKCR5t2qm4dp0tuv
RgthdldJt5W+mZaKiNGEbQZ2Zfp0d4GsyJRAc7sVs636puDPJeGRmd9f/rJnZRTwjPt6TANZYM4L
Jg5X3ceLov1404MOk5ZK9ik2nbZrfGNbJK2HPk5eRtATHBsFCmm9cKNwUoW5Vtq9Un6AxzyEROWn
dW4+f1Y/VV/jauvQdnRjBCCt5iIyiivCPVvcIh2swJ7I3h+dAGnNl8c7dnVfsaFIbEc43GLgiKZI
Atli6udbrMhhoU3BX177Rq9KEBCS9tsQDZhHnr8Q/n01E1dYneJREni3ifsFdx8SeJvqCddZF9GY
7GwPW/RejD1pSut1HsSDUtW2faH9iVG6zOtu6ioh8OEvFrS1jo67V7tJw7vDQgXPIt7kAuA5jcoj
5ortEgVYsc0njgZjSmT8azxN+eJD82mVKuWS9Ds00xlkfBG5es0feSlDeB7DAjv73i39aGkEXyp1
vjdlT1TlKpagMw5ec6F+jNuPgl0Fa1kWUdyOOJknsq11dIL/ZMSzzphpbl/pYQZ3zNCVMList714
+Fiupv6hkuok6byHWqez7EoO85BZfbAACk7/BV0W85bfbbFd4d+ca3nus/sBfWWA/Ihf4rxu+UpK
pCP/AE8uxQvpukb3/qKHl+IKwb+ygPXTz4v8XNCRICayOqjJprk8XzaCu9oUG3SXeDmZV+4OBt3R
d9AtEocg6lOY6CfqnMsnxbA+bVW2nszBbar1tFOKtWNLVbwY7TzioiLv0pnzaqT5iA0FTZcVKs99
KBNotHhhD4KMnHjzNjM7nuwROtOfBx2Tj/tZgqfmnO31+S6iKeg805JPkM7SNWE/3adQfvFjUjzC
B+oRWNlPi7EvrNiFVplJLkcxXMoR7Fvl6aJH/n64o6yDgDMcUKUZnWl1iHO6b+gIVscKtVsQ+NIS
fCjkLkqvCJsskg/Sv5KzKbW0N/I+8qcI58LbobkI3CK4c8Z4gZ0pRDoSanUWBdYGEKiZO79R15jk
RRP5bReysKmwqoMZ0p0Or9bzGV7gpqSwwSHgb9vpYvM2sBFwNTWltYepclCsc7c29g8hAQNttx/X
dSs5kjOSRN1Z6dFZrK9wNq/qINwm0IsLeQiQG6lGw+LNgDXq/9gbZIj8n3cai1jgTkvnesBGa4uj
Yk4SXSV1kleJCTcEGSbP7Ctk9oVisKQs473TLIilUF5pbMY3XzHJFwB78R2eWtQdyIia3XxY5y84
kMQNcdusyGNovwVzxS7oOyC9zKpCo+o0MDJ6pJeUDGyO4ZfDMDVRThf5oX25fdWhzL2bs3XLqtFi
EeE2GO77RnZRLhsJXqtXnERBs8lrPKAZpu2cohYTSYqbh3B8vuSH0KryucghfE/14izye9PYkv9f
kD08GnLOnya2zfgWUCviDcO5GhS64E96ZCsqQhZwuQT90zOwKErWVpcjw4gJp3Gs+I5K5dG7Kji7
uHKwPj2AnzupnMl54pTT1/7mpd9wug0RGoFzv37+fTKfeyWnFe/dFlkByXvv+t/zACct9cBYWz3p
chf9KV2g1B6tTAqP8xsPCCSC92Lx2pYSRM6uUqDHXyWB7h2MtlJEs+KrdQzXm8a91DNMGXTHbZp3
DdtiAxSeD+PhYICvDLEBmZjJPPaSHb8ETXLX69hQlwNharptWLOxb+nzP66DyGgWtO+umVKKg8Bw
Wf33460ajdMNwVAH8e7P8qJ1+XRxH1CCLbdJZ6ldJzdDG5cqwzN26cofM2bIM9ud8LIKIwjjKhUx
wT/XxMob/vdGf5F1sUW/+oBN8AUKyx7eVd7E1k2K0hwhCDVPx9fhS3UFJiTDg40AGkXl50PNfkGG
5tpoX1jDwet0sHb5TPGT1f0rNwfp60qIk0aZ9e3za4sh9xHuSO8q0qBIF6DXQsZj2Ht2wOqlfe3+
JLKTTbohD+R1Bbru/P+MBOcukt3yjugo7tRx9jOkecylV/Hw7dAQGePcjrnRZcRrz6xf7qdOHdRh
rFZY077yqPAoCb3i22qgYr1w+lDBBkYxe7m4XBNSKRWtpIA/ajWvhJygm2bDiSUZQJp6ROtTyxJe
AwRC4Fuy1ggsXyapaAHHVSwUEdRJWE+agQtXznBu1R5j3mQq4CGeirnlO+y2okaBjPTqelXY3Ix7
mphAukUL/WvSrY6lkDmVG3+KIJ78i34Fziz9wQlqgsooRVe+hdVPFNRUWBaBvx8C5GqPk5SaOMBz
J1s4Np90jygx6L/M1X2Tjy54cdvIxvU+FQStdcgie31YmmgSHJMkJJ97bwUuJNjH5cOT0ToarjpU
yzuFkvbb1pFPj4VzszJuih4kHpbbsGidUOx/9lJdxKC18qnjYwWPs5kyfxgIgT91ROBF9ecuHkIu
Gx86z4Szc2N9eQKMHBu2qRkpmqSu/miFFba6CxONlZ/w+igWLnQxGpQbIgATvM03t7ogtscR2A9y
x48u+OsWuDSE84utyYEW5t3dUcJfsUJY3CGu+1JkUe4FB7nYWXYCz4mtJ5xqfhvKXbaVtzHHsS5p
dOF5QLD768pDcoEv6j0gwOz/m3YCkPkQsKLm4JHfjl3GatbBmwHDh5d8cDzqZ6JvPyjsrz95Ndau
3qrzwAIVQUnx0gfvTqwn73n8dW/+8o8dO3J8g2uteOb7yXqMRkai1xMHWXSs13h5CLaw4vAQq93g
62aLg0YVnJKSBtvUQ+ALoUDmOEbM/d85l1BtrjyhXM9rb0QS5TFSA0wrXZ4KCI7cQC9iaRwtXHwG
8aBG+lguQ1MmVF4P+ccZuK04NZu9XwyCO8dyPLWqvy3/DV5ZqtInFNZWSfTiO/tO+u2izvk+YG4f
OdJ7LaNEc6mAnX0wVoKKFx33y3WWD3CYdTPiS0uqJxl65nyG8BcOOAuO7/RMwgNrmYfdxe8h/sWu
RgZTB4CXsMxvScPlDhVapx2LrbzxDgKkgEPp+M+LQmcBLc6/RjiH50PI0Qrz09hDIWjbkkCDbQcD
FQD52yEVz55qG+1XmzN3w5zHS7Q4h0wvS3h4NFfcY5Ywmh+h8xRaxFtnx0/xKRv5wVXTZDw1kbpz
Ral+UM+JwhN5HtsWt1wz2Y0AH8iXJpaOT08MqTUSWzaUWc1OvW9LL/Rd0UrYc2hCFllhiPHK1z73
jwn4VZydSQTkM7Bc8Qys56oRKPLxaXGb8S9V+HM9uhxV85CLXYDhfL2x7ZQUru9yMk+zgbMkj82s
4UNiJ0xjMicosNd9CidBUQyv37vqwpRCQpS1yWRBm+/bcn1+YBHPSn1DBss7K+KLQmQzK37abVDn
sZWYIPMz+1bmdssr9Ljr4dJ5KdYxUpEY87LF678LTt6Suep3CQkcVxXy/8Ss/9n6iKKWbo4wC6/p
1vySFrqA/uNgSIVn1UojVle0umC8Y37VTcpvvKcDO5VgSVddWCZQbMeZmNMAPhGAEQMI6nUUqbcb
PkLWDFykqLgs2cd8kxG9khRUVssYXOmh+7iW7EbPGPdi/5Q7gNgegyp1sOambJZlOHDY1xsxxY8l
nfaFSQflUSnKRZhS3mZ5BM6vzjYy3KU3sIMjx7nR3Eo265w4Ojfrtjwf3R606Lad1uwF60i6eib8
CFBhQFhczaqBxZyrEb81jzjBbqInagagcs/TiKR9dx83vyZHk8xw9zxKBVwzRrjsmKv6zckwCjH4
SsaMPPha/CaJEIpdIWABYazVp4eXKXHcjzqtWcoS0Ur6aYU+uGp18+vhXowbnHQyBraN0TdGitVN
2dLcxz4U7Mb81+p+vnxgY01TJNAL+cX1FcBTC2MnhYUTiDn7xN8NndelyLdLetP54srshtBQS8k1
Ssf+PdL6Jlc6VeTMOtVnoc99A9tn/W8bfxpvpTE2MOPJXm/bCTlrr36jtdv7PgQkyXHLW5G364lj
E0CfTPdaWzbbYDugrS/ntvUcf3/n3F3QE7+pfDO2/GhlOeE58hV2+ggTbwhmjaDfDpR/6gSRqDAX
ydpqHN7ldbzID8O3OnzvZG2qFc1izhIywJwknB17AzQAx/vSVcXSCYPa9JertYWOILnAgSa+cKd6
Lxvo7p1ziwrBq50gqjuAhC6QMHubBL1KEEyw27X8bCxuqhX87DbHvpcPr4IQ6U+3ylX43tOsKiCL
qdfoihfqcDbaHXx0/ln6vgULvghh6mZXkOhCb5958ICs9rtZKLl785GmjeMJTUKdtKxEwECelUqU
4dYyyiJ4fbDKeFIv5ShfdaZM5OsDZ1+fTzVXyiAMBt7Jx1NQcqS+GtGz3QJlFDmGHaSsr15XkppO
VN8o/I3eFqlRrpjYAvRfFz7lpux82oyJyx6TWOA3JfT7/so1+9qEKTmLBhtlP7Fv/irGgUJlcUXT
xFeVK78XnqFmHGWSDn0Qfum/UP3WD8Q+McTdtoT85fCpEwUqqHgSq9BjU/rzTcAA6kYQrthCK+Lb
P6D1/zX5zeLuAs/2ts8mG+GSaG2fJjZSftIhky77OU1d5NsT/xSyi62vWvGQiAgK9f8FvlzW+i8D
4vme3WU1yKSdJjmt5WEds6QqII2sVfpCeaTjQui3Hn5Y6uQfo1yXywEPDOy+Cu6lPsK84d4CiCNt
V7l8TJEct7OEQNYMutR8o8ToyxhJ/ftlHQ53M6BfCFRX/O7vZ1xRGQbpyjD9w6HGmGlSYe8X9kCi
u4XztfpaVxKfHv8x91MAet+d0CxJs9rYxvmoumKcfyco87DBuOu/XWWv00pf2e0Of/hrB7Ankani
+9EGMHFyljHV0lFq0r6u3ber/Nf1iKm9njm6zNnYX76noJlKjwgFCs9vO5ivO7rrn9Lg+tZYnJaf
z14RfHtE0UdEpeLSpRuNH5kohNI9YccjUjICC+JnOCLJ6E/Wt+fV3wL6Ng53lgR7PUCV7O47VmA6
T7vLMiJ8TXneeg3Q2R9Y3slM3oGxiAB/59QMR+niLN+Y2cG/fXF3yNgc1EzPLDshROklVxX09lya
rgo02Qjm5my7QmbAiWKT20MY0bQZKPvqFJtc4E7g/8ldI6PrvXiR3HPivZkZBCz556cZRfIkSlvP
urO+967z0hBFgwoL9mEdnFT/eUZhxdlbo1VGp+LTp2tYy3GkV4qregu/fJ7TMpjbXmh8R93TTSit
8f+M693vNzFKFRtsN/SrvoUJWacqPUhy0iJwhgtr+TYy8nyOsmJMyqkDIN51uC7HtgMCsjTWFLiM
6XrQxoh5o5rtFThIYp3FgHclJ2UrG6fVUpXAL9FdWmZjENPXGjSwy2/zYs8uPEGUZelzzlr60lM6
LF10zYfsR78OH0fmJnnV1KzDD+rhzI5cQFX4f3LrnlqdtlmXehr8e6rEejjHONC5gJEoIrvu8JLk
TeB0JzCZcY+Q40NRITFNWFwLgiM4oBn/NJhd3UyAlEL8j7KRanPbH7dU0xzvfqZ5Oy37C1ZubKpy
SY2Nxg7mAGAuFyKnEDLTPsaXr9w+HaNs0uPunjvpU0zqbLtZnMOB7IjZPtvvRRbxcvcsqh1ezFCo
9qdJZvcZGQP/beJKDdSJ7vG0X9FOhf/gr+pi4E3bs2+8WwG2nXzorDBCDnfHmsHohoxL5gMaKz6V
roaBwuZDgI38J7ep1D8kEDIVZ3fNh2N2QRGB/EA5ugXI4wUQycc2B2J0aZtlJf5MHhG87h5vqAd/
o4dZpqqhvV8WMvnlqk8q5jo15cjNVUjDR+17+GeeZ0mVroarsmJ2OelrhEocNZVy5F/hxtva6Hl9
qQYvEABVzg/eRjxBKuC6EIGcjwuQ+4z16s+N44o9Ect3t/OryF/LSVl9/OZyg+nMgwlH4UItsmcD
bZANN+KHXv4HcN0oS989M1dIwCasbvzfapCz1g9F7HYgdm24jl+oy8VM/tkhqS7wL/xrCJndyQk8
ncIB0fLDpsapb6B5QtDu3kT3ZLQPKM3WB5lNzNDj1SOe6AVkRxaF6fAm5Y2Of/qwoh6QgHahMQwe
F7hoMCuKNptAKLR6OYUN51WEgzaoW5nvYrAeF0tdxDfCuEOzdBtq3EWQiRBaof4ni7Gsw4HfP/Xy
mpNSAE9Ad6mQvqrqKAEkXXEUfuOfG1LuxHcY1PKyXvGLVBq/5PDt7XYLL9OzZv3jBlYbAkqpUW3x
9d6JAqI5fnYew2CgUWQu8F8ppwbNX9cV2+zcQbHegEhG9nqj7MHVPSjNHMYjZKWU1MqzFpoAHVd2
qOvEmAHQrGXe35o++SQJbTXf3eEq1J6iZb2/s9jncuLmBVm7P/Pt8kUEAUaENv+fYbJyH6G5JOvT
/mhBBtb5O6H5BK9yjacokGpCSQgjSL9pAPNtsgGSrdir39g3ASveiw3xBsV23/qYynx8yhCZx4zd
ucs+W6IA0uKt2Is6Mrcp2R3+2M282LvvN8HOEz+diORXg9TG+o7TY1mGa+NZa/BnwD6HvtkHOZ9E
7CZkOkyFXAhBo9y17XuvS98gSoNrbcmc3oHnDLgE3z0px5qB0k0MHl8VfQePHEPzZo5IuSn9WNQe
Fb1lrBYsoRjxzaYkTENlfhNSCQiL1SR0AIIJFESS5VjWesYuMp861RjUh7p0L58qUcOQgPCkDrN/
2aARaH1so3V7Mwqs0cQ7o7cjZBVwgpvGNI6CJO3pvEOovqWSHXvoHH3/TiAb9cwn29A3H+JATA3J
Fz8cCg3hP5XRyE03Sl8X8NCq0pZeW2ndsgcW9EJRsVXbhNVbbOJrhM1vDLxyuvWmGbKv36Go6vS5
XpGIjitY0xTW3DhnOznEkDMf7Ap+ldWpPEuN6O/xS0hGfsvoHD32MexjNpB9Im7rIy1J8HkXv16e
EzGUP6/OZUgP3kQ80+R0OX385rIXKYQ4o2/zia8f/N5nlzOdlxWbLY4eWbOLQ6TS9PUpSkmKqvju
D+usrySAOjZ1G9VVK5bojjORWCjlxXWf7LNH4jJFtoaJx4Kmb2pt1OtG5mXw63UBQfojSuCf+UCi
VZkQMwI13WPN/47xD0yKT9eTb6OCq0w09jxOvq+bysNW/yapfvzrFjDW/Nf4fWudANARqKjB7Cc3
w16l8ramk1rC6DwhcCzog9KQFQpm6/qFl1Xw8iG8pu6Xa71NfWNhmHONd5dvwLqAjuEcfv2e2DSV
dU/pGn0dZObjn/P/OFRa5grlyH5acfdYFfnWKSIekmJAkJMi/H6src/JUFeYPxGIdu1gWpy3k4wf
F2R8wB7SXAP4q4kj9jzZfaebgN1+qb6lZzSms6ryfos2fP2lA88CayxnU5JsTvnYY1vNwlKltot/
HNfl6aZEyWepHcWgQbsMbRmfRTpKYzk+mlTBubiD2+Z+N2YX3D0YTPlCwx952N5DY6F85V8V7hia
hmntt15j/SIPoc/tY5GonqBBhwYEzc+dBylXZ/dpjLFRps1dQCqdphebQey//qKJpESNrF1zGe9S
qfwthf9Sm6SY7TBJjX1hpbUNbcBUU7GJnnlelLnF11xzrm8rgSdrBjCYTEuU9xtTjoOFRwY8UvFX
W4g6ll6fvzSS/v54SMo6lWn00tcoEp7okwt4OwVMq2NFf9x+vyvqP0Jeb3CKZC3xA7eeGIo8oVpJ
JHcAaAd4a+X4wtcijjE3FqeOCXSdRbbqKzgb6iCAa8TLLfNTlhRXkbdnwVWkHmt5X78HtM0gHIMh
GAzUZo97/w9DnwC7Yl4yGTKU1K53eCX6zqelmYqjYnVmSe9D5LA94nKWmZybhpDdCtT27vrFUBCk
bLZ8EDNvC+j2cPh9qDcQ9oZJAuSOgaaYZ7A8zszv68QWT5F6RD1cuQZg/eM1y379G53uI73M82Cr
JoezPendshsIUKunU0vK+SUajy+uDUHLgZHcb8SE+is2xkIlFCp92raM8vsBfTXED2VJNryWuMBb
ldFKrq/WRPvPGI+9CJh8n4mUQz7oEOa/JEdQ8XqYG4VQtS0q3XBO2j7nvxeSZkNBqT63L/bwfGKU
lXTol4ySmmwYautnghOMt/E2FvamwPxNqQjnLyupTtVjcTFsXH0WSJu9CpXLLdlE2OThTpNpRD8m
GMTdDjymSAXxcCieRmE90Q20GS0RI+96UChBl1qfqZFv5bwoV6FmLxbPsXxQCCNtW9F7YeAsmbd8
VZ/VBZOZdC7BZiy/hT9DlSEIJJjTjyjPk/YFrsgRcyib9W7s3mpw+spDLKwc04kfTZh4P/5bxDjv
qK0RKAXjgOPMAy5TqtKQ5yPC0YEE5dAXYPATFkeRjqy6N2OnPFalQbomGes64zqIKYWZ8ufXxIk/
THU4uRWJcEbFsXJdMkugjXHmD1OMfOvBsMa0zEjL5IUMQQDzgZqjxzZJCKtnI1M16iLqmGhS9vhi
/TGg2e2VbQyGfSUdURRPljKH94Wmqw67pUZbVwyZfGI+KVgq85g9Ywr5nvLoD76zr8RqtZgv2POA
G+O1cxjiF/ICeWJT68QBD0vkc1wLp3LTx4pd5nsG7XAYvKkaI8vo5Um3nvAlNldBd3j2Yyq+kbwP
RTc7fnk0bG0oX3jv/ETov3MkDlFhPbhqusWitwOo/1KyImxGppgeVyyeCWUmx/44biyd53renbLU
fGxEgobdygSrIVYlIqzNS0N4M4gi7L24gP63WtcmbLxFUxaZ0opdrFMu6gXgYUW7d453c+kRWNZ4
UrMPkMtjqDfmG3Mtq96tOITJBdT4x1QzKk570iA6jBqP6WNZuPNyycYt+cwAqKUecIm4IlbqULNG
rY3lM8t5S2Ud4NTO7JBdSCS9yRF0/zq+Sv681o8GkE5Pa/HAGSGPRYDUJPEVGq750mGwtVO2SnDL
1S7mdhw43YatZqB7JTxmoPBk1+Ep4iKdDRe01Njh1ZGEwziPApxI60l8bD0ChGqDZL6sEJbVtNhs
J7lyOCbE33N9YXiLuFdPwbR5T0rZ8VVm+vNsKyqL+SgihhttzcM0dIwl19C7wfxmzW4jgoVRiFiE
SJXozBc6hAZVsQJ83AIGesdqisRtmHpCZRil70TgrV9tQEyDU6BQ+csIdGCC7cntdNZQtgjkOgEj
F/XZrBSpxOO0TdfqgiDap3ZiH5vSwjzRAdwn1nHXmN/bRGbM73+0uy165wiCCyN466gyTRuWS5Pc
w0yJ1EbQsQoTFRBtDlejwhGiTJ2SlS6dO8xMw/DYwOSQ6Bl5M2WbGbuPregoodUtdzcXkT3Ge5Fy
dtV85MrW/YufzYss1kUlq+z2DyNL19XtyWOaiAf+ZNymwJ11HPYN9Eg1WZ6iLqVQjgx9/c/i04rQ
OBNAMIvnfNV8ULBw882S0tOAlHgPSttlyR3o6Clm/ChBv5iFYzDLbDukAgXngghY0kzWU2Mb9U7Z
WxX2RGZLZ/sTfiYF8ESbk50tMm5T4wkpWDv1CbjYzE+8/x7WWH2qf8qjMm4hhT4C2CEzw/QK5Aed
DXkdORULLjkFa8XeeHtKyL9TgSPcARFAzvarkv4sQzB6jbC8fZwxy5OYst3nJHVr7kkmV7j/ghZX
s53HW/txUitELc8GXJQGVWwMmnxzUYWpSz0fIP1RvanM49KugR81CGgcuz5LCgLNHqpIn5LUmU8i
LgzgVQCvNLSr/I1/cNLOw9QvSjN8ZwvgVBj35sDCG7U3Ylejn/b9NSLpELjKnK+McwJXUF7vLH5Y
ab5z9zE1OobMsP+5qZJeu4T4z2o/W8aUGpaiAKNXKHRbPinKvcwP+SY/FHB6JhfMgEJj1TgnFLH8
GHVEbnM0uhjx21I7T5SyCetM9geqmy28L1kOOAv2s3C6lubrNGj2v4OP7eqDc/urM7+yjJO+RHIY
WYowc+5Ggwo+ZcXLRhldVsIESbN8toflLqrr6/5wYwBRiZRPAPSQukXcJSHrvzu8g8AllvY+tqn5
jkB2z6tomRUAN762AuiZATm5rdoXRCdXuv5erfB1paqdKbYgA79LTkttdajfkGVdn9GpZ+dIvBzZ
XpR8FZWXMa89FnvZ0NDjIHU4r9jO0TellOY5qNnIepBvmwObl3kNyTtYmGl6BhgjVBoBYjNmaG5d
pAnNRREayApQ7hhLqccPn5576Sw74HNedaW8LggOqIsGjm61dpIP2N7+2qSSiT621BPaC2i7HksE
1n2xK7CLDJMpXWL2+QMLdahs23DrtlJzduS9ifG+OWvY8Abdr/OaR7zwKZTs/ap8tbN7tkPBiqLQ
1ujWlDfSSiby06NEHMkWBMl8tDRf8BP6W/2XRagJHR9a8y3+/mCAwyx8l9xgJyKtUQYaKnyD1duR
17OiKPNfqgWob2cevaDt2AeDp8z36jdEZBQb8ySrMaJtPUssbXQI+LPrxKAJ68qDTWFYpYPJDayp
9DDBFxtmytj8o7pvlM4ZIyrQhw/ssOoKc2GWkBJRxFMsWhyuMV3o+AhtnW+1m+Go5MGEjpcKJOzJ
KxB07ASvwzTsef8/g7OLxZnYw/OUEJGhSHDEkvXjIqdmD0k9SvaqIsRprolnE0cI4FvaW9YB/NWj
Bfemqd6lZa9ZE2/2z+6bkLxNXUkQRDSn2SVCKW306hKHBixLnNixMrZQ/Fy4frvR0jggVD3Rma6c
yWBWXKKdn1husauIng33KjDxQWcfUHqwcB8WR5EA2weHtep18VJfJ1IoEoEPE3RfJNXvLAvow4lE
vJ4Q14a0zftELjg0nKIGK6lsKXJMcgi5XgoUxXm78OVVeSPhTQ0N/3Ctzt/isbCRPayUdBDInPRH
4KYQePQ7mbdparAK2Tvt2QyDp+O/HKy2g8bZphMUTd2d7nZDh++GItPMyhoRi4bHyoYMsPJXTC1Z
AXZd9S8IDHtBlt+M7QcuzNphRmMVNcIWJ6Uyo9EcVXySid5EeS8uuyEvYgmxdpcX8VrgSCg+q5FS
7eCstrVxrgDxxTza+SPvCOGZ9Wtsfg+bIgNO+HvWKSJLM9sjUrEe/2LycXWxk2YaglJC8IokkgsI
euttkpIcWXkq7ul9dUHpYpr18vO6a/8450lgy2+8fpyumHfLjITdDxoO1F4d7YN4PXs7EC8qbtzS
bExf3Y9xhy/cWvrOHKqCJavkAA2stRxZpzYx7Fd5jG40p9MpDDV2Oe4JJ77hl/AHg9jgLf/gX4E6
QSAIzJiLR+V1sSLihdPDvYvK9WYNSRrZ/yBodx9lto499VIUalk3C43/75Nm4x503XMerg0BbVDx
RqdT67rGGkF1LqPPuvRF/QVFSkt6IbMVmuFVefNcELJ/6gPN8nlLshRRK7XyWxvKA++P7/rRvmip
J+SErFOrNodldEVr171q7iERhX2V8u23SItF/4Jmp3qomQuzjOFXdpPO3QXxb4VCQDnac2IJCjuE
cr0wMoZZFbXEjX4jiUU7rLFPXMPm6pMp2WSCAP40R4mRmcKeKp7iKdyRxQO50H9HFdGm81bTAOIV
eveENFUvcclRYhnLWHjZeTJzX0tXT9x6r+vJTdLMbo5FS9UtW7rR9oMiNwDrhA+l0/9T3KiIoY5L
NQ1e/Cduh3EzrYPLqltCvpknfrVQtJs4O8f9symWc0XBbg9IJhulL89X4SbW7+xSA2jYQpsLrsTj
MKjOdjdKjeLBILQ40tdyW13gen0rQIBGmMnl/8PKJqreA32TJM1CHewWsd6Y5YJpWyly3Dxm8nJR
btpbI68ATROfg9Y+SCpEfyzJhE7qLpEFMw7INQitnt8Qbs7ia2XWEpNJ+tCHZ2Mwp+dYfdtkPqC0
6D3oQznUyJtHVRpDmoMvhbI7GVNW9n5qeVEMilbtzMYBx4pSldsVPDUAtzdh0/hAO7G76e2dX/d1
iu0E51F+ZqOAOjHANP2R1rc4uczNVWqRd/BeAQWSdIiPBc3oDuuDWndwkE7lpCPQUMdGOevP2czk
cGz6XK7/9TTpi0xxb96eynfM9MQwSqj9ynKQMvNFPvwW336Wp2iR74PUssazg1UtC/bxJAnz71mh
wmk51A2c3plA0tCXNW1UCbXbQg2BgkxBdTUNDD1kHWDWR/oFGQ6NP++iqd0XNOutfLwlu7WHk1h/
2hhBHu5TMxbtOdqqZ5yKDCgt6fOxLhgwMjroFcl20jdT/7yfGtXHbyFX8fkM42pN8YWYy3zgRH5e
80zmNuJSDj+0qgCvkP5QpzZW+1nWrtTV4QY03gArpopiGK7xwuLsOWrM5EMrL5B5CjFbP35R6laL
Mlw6mNuObLNpUtazDsMrr1BF6ZpKhsQUHVKhNQfzBZ6/87BOxvFoYcVETCgNyAFPquUAtn0OJE6X
Hme+qYrZjrQqBZg9ABzvlCYDqMNYTjHyuzdmlyeIsjKHccKx8YOWjN3TV3z+vqtAQi005SMj7Hac
KvOFRw8PvId8f5j6KNzy7IEdPyQ/OM/1qf8WKujsTr+uUkmhk8Nh3ad7R19Uwgx1ZEe2EmVqGChP
dzIcV5d+Hv0Q1P0JLChLvNWiWeWY5Ibl6WrxwNT/rgbIVjaBDlTPBTMi1vCoU+DWLVrqPzB4hfj5
se8ISvKfTgdgHI2j9xU7AYY/bPuOGF+3HdQmINPPOeqQv+az1YFwjGhRb1ys9SVPQNU1eqOiZD9i
PQ5PaJq+FVnqYIjL9xYUlnETZ/90EeAbimnT75cMVnVqi+zQ/+wj6oaqEsqCQRn09kk5rwHeMZAC
vokPSJrVXK2tGiUBSf0P4DagDC3nXA2xDQe3IbSYCS1xx7uFhhNUkmtudKR108lFJ2FtcUP3IujV
2HfMgMlpP/LCniGFB6tfikL9Aq2gqITYHxU/pBTtsH+DEwGar2pHC3y9MHfGpfx74rsdPEbE9Q3r
6WwVQ11ZC3ELfYCARS+lOO1c/PITFcVR/PRhMoJajORwtoMapVBg7SAd1PHOl5j/PI2JYNGozvia
fBDKMusA9GQDZ7iPWo3sYhOtG0y/SKdwCWt5Osh0yegjr9tdoyr/2LShUsuzIlMMBiNMkHeVFXoJ
4ro+sz3HcLvTXke7USt0K7pjOSL3/q0iiiFbaLIsBV/t/i/vaoY3qCA559TELIrfjJM5+g7re+em
kxG4pCiQkkhrkJjESwUyBcijDF0svrwl84EmIpL6fld9Q2jUnk7oJDCNnhkKa9sJGspi7lVZm2OC
xraupaoPWP+R4A1hhAIr2yNAVGlhCSWR3bV0qyv6EcSYJRp9btdF/kY/cFgSMic5BB3wM6oBUyXI
38IQ0CNYrJzixFKHm82pbTXGzgE/sK8+ji73V0/9U+ozlQGYSNFOnKw09X2zF1v0XjVgHtYRrezg
kW9yniNgrcf1HTfgl3by8WJgve8NNmqDNi5534w5/X9ngOC3lDRStt8BaQXCSB9hzmQECVQHSfAi
8yVWY5oaW9SCPl00wGihEVTm1MulxKv3ZssmMMCGVG+6f9KCwUvLGXmE8embI3UIwpvlPitvz/U5
0iSHSl4GocaR8BIZvhvRdoVjUPJF7sjj5Ish0KBiFUCM3qoguyjILTaJNKXrppq5Pc6W4C9Jm05e
Y9gGWFHP3+jcXTtyEi9TQcHE0xeByL+DBIPxgDs/xohDrjzUAtOZLGF7uykaQ3LTuXO56ppyXL2W
dcEbTU795DIJicVRhHxZoF2XOc7RmOmL/g8hzQUpaPCbXsgKgxMZixtUji7hfypGO8msvKsvJRk1
jHY/0hiRe42RK2U02I89hIGFj570+83XDPnoVOZ+qiGVouhe2Oqu/SL6nYymBZbmKm8202O1R5W7
PUjFceLMELbdT5wNIf0mRG1I3EnCmCIfs5s5jX3vuSXSJq7HAhf32CN+2mBzSxI5K3+1FdlptFWl
u3TRN/3QzG0Hinegw2mac0sSLaWoHpn4eEcYxxGqCm4h1XNDNCTpY2m4NyXgcNTvccA0gdW2eGJi
54HY8GbDBRxaQ+d6MZX6hXzPx4B0kXA6K/yF8nRf60W4T4tWlzvEyJXz5oxufceUO2yVd9SnYiDF
JeuF2lR5uLGP7RGDInwT46FpFhJLHNK4SEPILx/f2viRQhAu1n/VKS4IPhdVOUB8zQaYRFBEPydl
suGMsp8vKRXdnQGCI3jjJDOkqf0pNMO7NGxwywmMqBtdqlIv361tRjVhlmFzBVtMW050ijuu+BDv
btvfi+W2xfVFdHBNzaH9gUeVeL4U6r9d8doAs4FckPUnTFqLAmZp0hwsNc0guUTi93nSod28D1ch
TWOvAueVW7UQ81Q9sRP61q0Z4nojTnKogY+VqkhDQzRQvKrTyuzp4+7HwQukvMm9SVJYlAzhYlfx
uj9Etc/qPImEIIbaIUCIHJG/0ynsLD+t2/Wcqs/TGQefFMk6YPBPkds0n+yanzsqLXM9x8nhEJbX
QNOae6A1qIMAzDsA6NegrsaAL20cqul7g/XiLPx9clRPuHeM0Ady83hgDI3kXjJldhr9H2NwU+xl
OezOWDAzVtLpvFSwenVnWhNeuCQYn8Cd7aq6jE43cVl2Vw+I5VEBD0nKr3OU9QrRSalXGIdBkVUz
OfMsTQdX0RUANWLUfxsIsAm2AgY07WHfqMdQfepAD+6omK53fhscC53rkvrxD6MjVO9MwivsY78I
9HCdFsnjaFwSRp09KFLHoyEn6AKSxtvOKWTIK8MUcLcCfDChS5QogMh6PiirrvNXNzpey5ZHDk7O
AcDJbotMk2sCpmfz1FIqtReuwZnesRnGadLbCeElrl7ee0EBPayn6ZWmMIhInSHt5e2UrEjeBzwN
HMNdB2+3xjFQklfJGyoFfT1NNLPZZNkiuHa20wl9QlfTrYJ3AGkc01JIyyhqHNQ/xzev2X3LczUy
FwBct8gukpdyRScljjEYLNq9q+E5pzezKtCHb5H812zQzC3swZVwMlDIsvJPW5LSOTAEKUN1ax6S
yveyCVDAGqDKSJeg2o0HxH4Yv8FVITsi80bBbvbbXBx2wQHcShXzrjvFQCGqmYlFRbJbFSKWNa/S
dYA2YjBYSaZs+vGEbwRC06g/5jcLZvMs6AIwYDZdUwCS/Gj2VYVhk3JQXk0kF7fW1/m+YsX1KZht
PGWh1nDYC8TR8MwEQwqIJ+tqWDBNKjnqtT5W3mDw2HlWUlMr86uB4daFI4AOCnml0cCpbuqO0BXT
YsOQ/Tcw6ZujJM8Z8YRdyW7uu/NqJbxGSog9GnKOL2WugFlEM7rixM8tVfw4+Y0Z3dm/Ct15XRz2
EI8Yqj9gyiAI3lk/p6GQZ7eLJdJqLsk5iIiKJ3z46FNiVyUQ/jzk3hUPbEAFAB/jf+azuTNNZLDp
UCzlLGM5wPUm8HD2LoxIPU4tT6IQ5tukpMvjcwJ48FsDVZkV3w8LHhJV6ZAchyapEfU6HSjD2+AO
/vQBC0OJdHEHp05lyyJMANtau4NXYFxD1blzp/lWqnnIXmeLeW34Emk2xDCniPTVF9OTC9Iffw6i
dmPSI+Gz+AZTC6REOVf4OLwW+tD5iLLZZ/tC5EK8Ac5sHN19gv1IupP+NJEs+oFUaEcLJa5waWdB
rYc4VkudQBDpiW+Hw44Us13m2uspcJMFfruYvh4TMqdjB+JA0DwGzabqXXExbPshNXRQyF3SM8ne
rs5yFOBvl655HHczeHZcPcZR+wHe94zR4z1Hlyy/YncTF05+gVwlpvXqwHjwkBaccO9yExQl/kp2
YThMfpJHPD0EvInVT+ath1fAo9O6q3LoiSuNcvR93hGfzwmemKKsIHplX2U/FP+5x48S5ofduMp0
tEpjbY+UbBhUXlz77TMTNOduMDUSLPVNz66hJG+TAIW8SsbesDDA8A9DNGsLAGXlJSoHKAwRN5Fq
DZSCD9IYt6IgjN6PfsBX+fC7Rpuf6Gw0DY6EEuPE3gsPw3rXKp66QV5U9R15Phz5/snmkENhWsv1
H7OEe4OlphZlZtA57W5ahRVIaqIy1tjkoCnXLSGYTgMNB6FT5r2Z1FzSTPQWH2xU+WE8q+2E1gEv
cQ+4Tmqu5msZYrls4JFX4n5fozcKCQuJ0BRienOPGcZXsgnm1NcMA4+YD6keepQ/aIWo5e5kFSb6
/7eXERfhjhHYogsc5hSwwNoadKwK+ugO31djh0zmXmbwKCNe9GZXlxsrWIeSK6JrdkCWM0m3bXXg
C59vKxqgBNcRHeh8YwUFLzac8liqlgpk/AViaCRwlutlI+8woKrS8NK8RMlabC4eIuj63BLAIyS+
o6s7tgW6Ilbxs4mZ3g6KCDzwmV0K4oqD/A8sVShYAcPW1Oq1MQomX5pLFrNGEpOK7GwvLYpg/+sT
EvISqn33Ry5JqksP0h324oiX6DeRbnZsZU7c3KNHwV1vnGNLrADybilbjVaGBaD8TnyH2vm/1ZMa
sB0JemgYpb2Ol3ZjRMaUHq3d7+ZnGuBk+uPZ8nCZGYMFyhbs2kXc1/WHcaL4W6lD+u5cXxTCuvLe
a7GWvf34lYW38WS82/S20OLtqfuWRndOW+1fTTl7l0Fpjkaf14A1bFweyx22aFTZapatadyR2q16
ibX3C5/49YOw7rCYIcrOZIapgGArse5NDjCpUgsbWd7s+08WAiNuAkMXtJwXtDPxUu7ZFgjiiKMC
vBJkX7QAsgiiqmjyIcIAYRCGmWqizsOIVVD0TiWrx5IpEqwSLzm4suZUouccyhW2GcmGKeGPdxBN
jIhBFg3UmFb9Lvmt8qxYukX15T+0gKrqnT3O4ZVBKwJT+qfp+Xtt+d53DT6AIpFmA9w9/BpT4sIu
lT87SVs4kKJRnsVwEJRrTm7+wPL/yuIA8/mgcebwtqogUisC+DWKLkWfUkn6e9XnPoT2FwfW/wzR
QdqCKJ1VWDCX8jFEN3eVmXRNnuf+D7pso3Ey5yZvPSBtrOgFUMh+jQFkNGeNDHUGrCUlAFq14/pT
Y3E2uB4R48OpboIIIibHbS4hKV9fkZXIlmWzp1csqINPR1BPx28Wz79XbNMwRXma0BK+93Q8YOG+
rvq7znvzlWBsJ6fvtJBFAzK1STlIdSYd9kJ3ZWRAyQglmgzEMmdzV8/WHLwJdAXwzYOx72tzDukI
AMrL4oY3zBF5dXXH7wX+pFMfomw97/Tx5ktOIP2xA2BNauGJG1CiN/lm1YF7oh/1SrV8PN1B6c+L
kFleGApkcZRz90dFZef10hP1rzZIy2MGdFO89mFsNdT/X+jdQtojPPOW7uALTBknOKDWNUfGK7kn
zXu1TpiIZ2dxXRjmc27LL3LH9xNfzGhCXJHkSRTYrIVWka9UG0yiNncH/JExeoeOWS1OBN8D6X9J
btjlMG7JBTum4Z+yu+29nxiCvBvxWmGwBOC1qT9p+HiZllPIbo1CuKTc0pvs3MvvLk9+Nsgh/d2F
C4FN4WZPiJcqcoDE2lxHFcn9GR1MN8uUd3nUrmPk2VqGv6coobjO7tbKN02ZY4IMymKVrHboa7DR
wPEGbCGiqw4gWuB6KTbbw3h7js0Ck9hOzxM1/Q6oC4nV0PodWbLozKGKF+tIkp4fwNetbVzvDw1f
sD2gVrLVhSNfKldEA3X+pfgfT1oTnzmI3QMpkVINUPhOH3jPkODnpRWcWMMjETB0PYAXdZQaEzmK
pQDL1QK0z2VYCe+pDpzxq6FWHwzL7tX7hg/QsxClVHen1wFRlspHxyFYmJmQ2dZFDDC3wwO35zGI
dSq0+uII7xVAVnmIYLACBn5QKmCGUxfVLU4d3rktJZpQIX/GRG9dzBs/c4OsMX/3zFBTdNTdrDig
N0RG3MZHxpD8M+CP9cneQ9ulXR1qGlzjBiDRMSeMIpC+gVHqKPDzUOfuLFxAdo6diYjWt2VVGsBk
Y/fndWTrLkRwISgHfzZl3MoLFotyBvO3/Ntr15w4LBI6XgmNaHq5uMemPuJGXBRfnpGgoyYKJTC+
ydM2j2BbU6uLcJ7D3/P1mRzYcMy5iE/P1ZsUH1Dvw33sQfof5bS1wFQKAMPjkChSB2qQ2hRNSNEI
SCA1cYLnKja/z6j8D8R1Tvs7rpEJnV7I+bKjTWQApCKsVFT8iBeZpVhS+Z3ia+FKPIoNFLoSU0cy
B7xbS8h/IcZJ8AESS832CbFbQRHYR/+393iOAGdohYvsWh2I+Mb7MvQyNZI/qmPGmo48vMijbhFW
zFSk44oqBCsqUI7tI6O9fDeVpBVT3v1VscL1kKslUVFtN2vBZzZT5nEPeGPwZDh6RsFMpOQePJM1
mmvVSKTFp8cKn+LIc+Zp3ZXE5G0Y33JBdMdeod9BkBmuMHn8SaPom3cOs/PRWc8iA/I2dl/pWS0D
3Re7QP6eyyFAqOjV4r3hxwf3QaD37a0abrgL/IG6Y7fuhQ/2rk+wJCZAtyU4m0Tg3flSPXWl1zNq
pZlG5D3wLdLMqbBqQxk7qaVu9ko3RMmM8VsWw3xTVaZn7epibtRDCaoz37zvLGWIKDR+3gOBndYH
IQ1j6XqkcLw6htMWqU5WqKr38ppQoFzeQdptaJyrDALEPeE2IZYFkPultad6mTJ30R5GsQgoWGvo
HSLCBTxEGqrAx6yt7IOPkPmAlLUowX+Tn9xAWcv47w3g/n4lhm0qfv/NvmJ7/pMOtufuTiswRr99
kloaXH6uBiCdfwEEEBa5ycL5UNosjEVlc8RC8i2ltZTvhL7my5KNBhCd2+6dquZtUQJxecKHq0HH
MKK3XNi6yx/nlR+2NMhIcOUx92YhHK04griT/uaarcw9ZEUDpUVM7DLQYngyBq425SQ6qZEwlSOL
zwUg4RFtNAyDNLIl5W5Gtst6PE3e+/ZE/IE9sCe/s60QPuXaEuvNl5LbuhVY6vTCnCKTljHQqc48
5+Ln69vM//SPI8RRob+QoRWxtl22cx3RFrCIXHedQdTHt5/XyUhQw6I9Ng5i4GAFUwLXJ7j1ERDe
lZZMfv/oIEQ/XkITKNhRIV4ddvAWLQLCQaQQfr+JJy8NbQxmG2jM9VLZF2eaigjwHD8RUpu8IaZx
LFm7oji6mh5GTkzrG2Ym0Oj1WKmE47ACvQ5VDQlTDZ+K1hKMAJayHopq9MJQ2YYc+ndS9qPcdyPV
gH0xt8044MDMmSIYcGD+Jot2je7u/51D5Cxc/Ah7TqeVU6iu2IrCCQAHp+8ZCW1WSiHFaO4Nawo/
fAHE3N+B3kv/BBIPlY/CkSmREOHyzj7zRJ739OJUAuP8hpFCfUzUQkke5cZk2AgPCa14lnIDxs0v
G4HDfkHfwc/mGrsMGGdykm0mbeMf2FX9qzJaH6aV2vTCMkkv1R2hy0zC8BNCNWmq2iMQTE8zoOWj
+RMze8qEslBW1OlA6fzfT9LiTiRZjTsAFsjXJcAPpMDpRVB0cYgewHncMlx4ox5UZd1m4B/nMukm
9xkJdYpnTUP5sLF59skyqjS2sA/2IsgQBPq4xbjfwXX//WM57+QGGOzhHQDEwM6Dzr8LrTpfnEoW
zqLNw0cmJOjSTYQTcM44bJbioEZTnD8rE/1Jg6gwlWhfxK3O24D9IyhbAxcYKoG4X3xmRrGC3sSa
V0KKgzmm3MPZZrznmEVMeq8tSy8SYlMjyDnbh9OOHbFsSogWRvYEpbiBSKk9t31Vk5HrRDdcm2JN
8ALNKnqig6QNLhFFSqqlMrPFgQXUDe+UXaIvBzO1rHIe7iUSTaGilSWsgasA4lfU11PLEd921hcV
cm+uTH8DPhdAgabopJvlbs4kLSNEHMSdFBv1Byob714Dh+A4D7CXtAgbm1mV6nIRc8una3OY5dgW
L+IKvgQP8M7yUo0WrDOH6SbNf7mPiR0yMfOd62G7flx+8a7mvHAs7ND8eS1lYa0Mx2mzbe2aPVqn
yqdWvPzWypubRx1OziI7PnkmBmcMSNBr53bxra5EeQ/OBpFuDOis2AcJCxM7DZbUHqeLa701vIs9
BdBOk+CzRYqw/GBnpnMjrrQ7LBrIOXkia/nOgLclOhmkvhk0TtW/TTZu7fd7Onexe6fLtB0H5SJ9
aQ8EgdtNOLhm0nocSNFXCVy/kY0spkCPij1rv6T3eBo672hN6i3bxD0+GE7NwT+oRQY9kFm0TYX9
cqIVRreFCGNW4eNt3MoA3dbeCX5ieAWYvzdCeZKSP0roHN+XC5Bc8sUF7iYSXTgZfMuSILvvUuAI
fdkmYVAhHaaXZ5zeyQ4JkQpFo1AhtvCTPmjeG887Dn3Y2LZxcv8CqdEnKOsX64aU/fApL3OlF8Vk
m8EXHpT5Z9ZW3hvTmBM4MD2UfyYkONSd7PU/MsZn4KOr08xTi7ub/emNHGzIEntKC11AxDazNoTX
fmvMXBnN/qxojt1mloOGa+okiOI80kZCmTbgnlg0mnQEO0Anw4g5JZbCzPFulWLXWp1ULJuI8a8h
vSNJUAVwQ6icrfES5bbWykSqY+bjVetnGubGUxdXWXQyAKY3qkkt5B6FX5TMMDhoVgnT8KbygwHQ
J+gmGJZhEc5e64WwGXSduTrYhDPHjeWgTZb7yXJ6k/XeEPpTP2vKrVPYSId1ImJqYSn7t7RB2xTi
LmYLIuZqhjF28auyKK+2vQwXpg4UbuS4LQOmy7Te/2imttpiKuKh6pnwhADa5AClH1qcGHTvMxIO
OgsvEzQc22h6mSJ17u4liQ9olA3c/jslo2Yn07jo+nJQ8lU3DRZR2me4HzYSfSHkg+Nqb7dEGOFm
n+R3N6Aghm56ccJdES9C1CWIsZqdCTbqIeB5BLVPfgNTqRvtUjvOxSVfHSPW2idK3OovtppuR5+U
ux6zm1aaKqEuI5EeSgk3wHrDTQvNh8d92EGUgxX2xpab5i/9iHEmwsl4j/BPwxQxh48pSLnwBHPr
TSh+Cqt3bfCykErR8SwcxYKSGeH3039+2n6fnBUkP1x0fZfKR4xjjBV2i7mo9EMOS1zUU7ywBcjO
bogkK509q8afohYVenSAubDs2zxaxozBhX274nBbeu8u+LtqecOjMfU8qszoXMVR+Az0YTsk0tRD
zvS0XgpMDr/uIgqjBfjW5o5KpDb6edxLn64BGCpj9QfOU0KZZk6uTB/AYOgwFieKIl2eDXsPksuR
wgLULB9qgxgs3/fO9U19HtJqwXvhHy4FamlfKkmkK9BCgSoBHiCngb8zMWjTU41/WpM3GvHF1TTk
AqPF/Dg3j0rtN5b+mnhm6IC5eQ9eiESa08x2piSY1RWY+wMCjQO4FMfcp+ptgsGdVJs4m7BohZJw
iK25WH9KTxCxolzRc2gxrZjZPp2P8alxHhYWkDA+nUFd9rOizt+VWhDtW0fkpv/VV0srldwbcbpa
T4vkjKm2AtvdIrcFUwSnsHoprsDHcCEuJIfs7euA9Tle9VTiCaYYV4UdKakCDwkOTK++Ks9ZuTGF
F/VmY0VFKk7hAlHdrV09NAC1KuRzRQA+96QClml8Kq3rWBKhR4ejkWGJyziyrpfCklpSW0Ii/cig
awZkAy/jOxo6uT4Alqa+5ffXAnCqFnKqz6RjDMWwFiv0P0c62y1BxNMRp5pvSBnQlK4324bZcXop
J0dMgv8scIP5psCWRiAFElc9mvMdH3RMHWvusQo1ki+mEV9dL3BgpGJeKzmcel7U/UMRcDhbB/bQ
glq8gcS8hdbFQqPnKkfaG0Xz64/rwhZv01zmPUV5x3M9qBwJr8mEzbf79PLkui+nQM3Uc03JyzXV
OH3M+G1ilNqcUNWGFBnpv0aFtyu9Oi4+hMqFdh9tFJdm9zHigMZu/vEzO3CLnEBUIZdeBVB+5K5R
xTVIqFC+Bp5RzQ7ys415hfx4MiA934atyhlrHBaiqpS1nrSbSTZUcFB8yOwx0+Ili2ynGIryFOTB
mGLUExPM61/ypevQ2XvhS8D0WJagqGM89/iloTfQxdXk/RtjOwd8o60RTdoebkdVSPJl5f5Y+i0Q
4C3cNPO+XU/xQyi1fgOckqs2NZtDBHjc4JTy466wvVlb8HZrdkACKjUK2gMQxF5JiGw9cdsxs8JZ
8i9m1SOQFMVTVG15NZG5CF7vrjO4PJD+Xs2/kcQrEWL6wnQA/n1s3f9mtStcmtJdPVHfUSmhtZcU
mYjS8OlcEis8MKY4TelYDJBxCb8nmS7Rois8wdbT0+Fy
`protect end_protected
