-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LSk/dKoDoh60ztd2tc5+LJrYZH4Vhx82kn6SCwUTVhL+g4gWWrWPxk72g3FvKzw7zX33o33EKxv2
YCbioE4+Wsw314AW4ac4Ml6s5lQuuZ2PKN/qvK/DcVBmKXznBP9r42bDuXruiZBZtkAKv+mMaPQS
aqqXRmxYJQHUc6eZIMVioKg1BxwuMVw/xsmItWBWG+J6w+RenT9ToiHzqZE1TU76y4omWHCDji60
AC32jfcGDDndRb6rEfZsorouFuq4AqLI9DlwVp63dms7VsnfsAO0kaNL96mx7GzWcvHbkqfg348F
gmDSl2vVOdDednEQuJ1ny/ADqQ3ZxOwQItE1fA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4528)
`protect data_block
WjrjJtqGF/eO0hcQvv/1Fv/QIJaDHSdyxq4+NLSMKbJr3GDwvS4pX4QRkd7XymrWBxLEpImB5YQn
0ctZfwcmyNcFRDQEmfHc90IjLtS/bn36abK+7OWu1rehfEZhMMtCG1aN0fq7q+7+gCMG/a3Nc8a5
XTQ614dmHAJLGXNn8CPdhWvfXr4CO/uVdKlQ4tl6zxlScYhWREFu6HUAdk0NUR1t8+nnq8RCSUFI
moTlRwJJ0uuWl0iJcG8gge8BITOvL1zICaqh0INQOrEqV3bNAe32/dOarXq8Bf5JX48lRmAol/EX
pjH4dVLEYIGYa15FuTpA3OfnodrmmvhJ1FP3nzntixdafZy9SsKaRirMBLnPb5Zzq8zbJ3HBhxb0
vVmPg6Ri9M3F3YBXqAOv99KOp7LSJb9GiM6XGjlu4ZYmprnagWeP2iAM5U/KUncwjhqm+p3gMXeW
u+hZpqaraGksKBK+31O6LhclciYM1bQivvmMpcZ8Yas5AsZOmX172yn/V4lbcWHSr5MefYGCxXTT
XqD4FLqp90Xt4+B6U/MLNIONIdOvf36ZbmKz5JWmGh5dS6pJviuNttGz+xjdijvzk5cRo529DKHq
y2QgbIKqds0AuPeJWELlPyKcHLADJYEcN4DpaNa3fXw+Lfz6A0EW5KgT2x2Bht2+aTtlFu1LB3cc
B+wPXl+pzp9hsFsUabcoy+7/j5thVtfvNOz4xscPDct0fquseObuoAtaHrAQ3ojhpug0t/Oni1Rh
EZO4QnYzNfpC4tWbP4cAnOH9avYcOhtFvEk+bbxylP45sVyaell1gN1jyyII63cRP4BNoEF+SDsU
z2ePhUyuqNYsVZbQZXw8Xca1nvwJ+NWz5HzSoa8VpCxXKDn/m3JbMHSOUCKPNbbyQSf6ORAjzBIr
21zzrcjXxSppGX6moavO74YP/nYALq+tBz+LByPtqWL/Yul7F99SfCvyMXTKyUpHCvXIvx4GgY7J
2cR6FjYhhvDcPjSMJkUF5iCwfoLJ7sTEtGsiiVBFJ+KtqYjHpSxX5u3kYKcSjUK5e15ADeeTiERM
QCNEWUeX+2Vb+1r0d/sU/1RdO+RIttJNmUoBCULx2gz9ivDlOSzJfqmJK7OmIDaWA1ayQJWcQiA5
WDiTP4PneXhH23Nxcso2Pmhnjv4kG21w+Q8T6W4OPE7UUKPC/8lQxaDDSSc0dETcr5+Buy5Kcyo7
aJ893R8lqpfHx7bIOGeTEJ31I/9T3Rjgm4tTPylqFr5ONZIXIQK2lG7GPeSiT7m0pY5U2P29z6/l
aAIG42DyCLJrnHRo3qp30JhLcF1I+CPOsRmZRf6KA1rnh4DIbljNrIbnW2YHs8SessTxd7lYFiaE
9m3SydQz4ysKbSM87Ddyjyijx/mVHsGlb5a0TN7BYKSneKdCCB++WTdtAbubuoHJYnofqUmIepIx
igT/bz7BS7Tvu5ONvD6c1hm751TYjV348U2H5FjfJhcm4VzSBH+3Oakz2imImUwS8kxdAvVItQ9H
lu7LilttXxxA2ZIIjnMMeT/b1h2FWNr6oHN6BBkrSJf9b0XFLk5OwQGos3hrHR0kgqvZbtLcJLPh
7wuPyRPVKdqnByixFBqHq/NRCnDMKJaw7emKJeGkuCCL3kyPNH0z9FDkZL3bVE1wjblQanLkuh1h
RltvxOBz5BbGaudXOTODzjxHoj8eOGMZE5vVZJoLI1QyG2S+qGi9pnW66UbvHiBhOriwzzVvqvBr
P1DPwhdrpl+tZTl3yvqF8YqBxAe2PqJArXwAxAjvqN8IvXEoQWNN4/hbq5/bZhkWuP+DUPfU9++6
KIK2rmZItwWYMWJCHBpgdlm1pDDZ+YMiqAoFnwGQS9h43eCnbD9bfcbBt5R3gFm41UCi+A64vEDQ
GvtEzojWbFeJBr6+OTzCsZZNuXFmMFtjQmrsLoH2Wz3ID5z2uwwMHainkyY9IxfqTByH95LMjF1t
JsWFrgwLwOF77YEkC0yOYdffl8Xh6gS41KHQLpDqVGDiJCHU58y8Klx+urkyzreabk/CqeRYMLRd
mnyHdJXUSlpls5TAX7AkVadOSsnITQekPujWI2W6fRAqL2mhhgPuEBmpLB+aqUaH3Ky/Av+ffogh
kXf1mdjSmV43Cqs+4eGh28vStv6v+kextae1nmsjmr4ZZClHbuo446xtOzZViLZJzyxBcYsUmtSJ
+sk51ggxwlXLObIUqZElysCDiID6hZGvM88gMWyvnaEFpJQL3mtekWgFsTrYRW/1CkqIM1HUplvq
/gKg+drucR7Ap0kMSXjz9ibBVi90tU38YhsDVwrb+CRsQM3hQsI4Jxt4YE7xNu6no7K2LZKj93Cn
/f8HHX42BRePduDp9KLfDToyo6ZPQvh8XqnIuhmrTN47s87AMeuEdTmrlrSYLR4LteY/inyq6ls5
n9Y8n6TNzfseKk1uRAUeXBqDNidG9xu+1wkTxYvqWG9UlVgDFGcyDgz8H5+J4fE82h6Qy+pQuMtE
vcwmFnSiKRCcqMQBQX3TsPPAR3skogfoMGL20n6cf04h64zKEpkrycbB20MVKCrIRDnwliqdGeQ6
1uKNZW8br9y6Ckk/Jop0g0oGSKlLJ2vHp3+cOeaXX00nj/ZAj9HysTorRIOYVRxc0xP00VncXScz
f0eBdzgtNIO46wZoDOiLwJdKc3PW1O5pki99qAxsdu/SavUNTZkBcuM0LsNvHUDeD8Att+eZL2F8
tA1jl5O8DFlH11xM3LG8VDG9Mm6cHM+yIaDl7BQZZ5KsR+ze9c/cK7UAAw+6WqvpZuvgsnlCVc2t
CMlNaTR3tlhw/Dyd5tfr7O8FYZ6teXtZuqE7UmB1Gf4a1xI20xB1uYXqVTD9PTDqhKvk0Y5JSz6u
C2IoJ9SEK6N1923ERExt5pmpqoAjarMQzRzEmvLw01FtDIG8JH583O3LOmNFAOPZ/s1wEAPByd8k
W5XG1zPeisZIAmWkVz0wl/XWRBT8BGlp1UXqKP3vFgVH/RpJ2Ju6lDlKzbcnNd3Eh1PvZyn915Uc
OVr08cu/f6tpGCS9KZmpG9i6iVCcaS+9QZQSi/bIPNOIEIH+bkyXP/Mg8vd6ok3G3a9N5j0GDZLS
2xut7/fBdP8ZTEhmK7aYwo6IkHcSR/I2LPPYWGFT7pgLGP6EHt72KxR45mjcxIa4Wx5rSMRvOkij
TdXijuSJpem2FyrFdAE9rAGUOoqoyJMjvDJKRHK1WfU8j2/ehv5BZT6plXAEuFq8JMW1fpnOrzBS
FhM7NuJbB8cNBm2oKQea6zOgI0WBz6nwBpb8lRfsn4Q83yIol6FbGRYMmHQcLetqPMSKgoEbKmI/
48ICbCIvVV/pJO1+UIv5g3vcx0XtpqsEsdS+aVefWIOvfWmx79fNF8tXwLN0pj0ct/i+hddKtRei
sAQJ4chFh3VIbHcofoGKDNbovYYt/4HpoEoAEabaBaokVCmhUE9g7frAQlv5uZ9bg1iw9BIrag7N
9r4fvQdzGQ27BipC2LX3rT1DiMaRVSQRqnZnlKMvccJUbqMdT2NR2R8Ca9sE1RxYGQ085VfzNJ16
XohYq5SmguvGk24JMfljkhk6fNaD+oVgofsui4LyZlxROj2L91HnC72e/5OItfGdaKxhGQQcbRbU
6csf4agS4xHx/qw/zV2IXH21aX2tvVjo4GITV2NMXz8pTCdxDeNs0xgoEf3xoCtwsVhyXkljDSAT
/GscyMr2YPEJ/XliThbBuLFSQ5TgG/Wm17E5KZc0/dzpgseW72IOSXOkKT+7GOCG8dUrANKJN53Y
gbyhL5hDNPqKyMIFvAAhOEtN2uJUID6X96NnsdlMMNXT4KFxbQtAnCtmn9dNdSZB5FV6B1050KWN
c6WaT36RtMo5ifGKD6Qmkk/G9oN/NacVEQzfZYu6ayGzOL0sDNzB+tT2mQSgWVjkpHtOdir/FzIw
Uo8Bw+caBmsjKqW2tDBIIp3b+4X+WLwfGV0R5NoR7XaJ6ZHj6+EAzH/LzRAIWxAmQBMP11+tS9Ef
1TiKCsNluMou/3piYtZVNfRx6i1p3NlCbDPIcrw9UtDzER9Q6OH1TWnYwVyuzY6JoD7y4vcl0A6o
QP0Z5Y/gP2Gx3UktVlwzVmQKPxBTXduEfXWJbizJCIpxBtiWa/Rq4spUnlENwpfWSQNnwrNL1SiU
cC/iswbMzuqh9LicY4cjwR5vafoVELCjp6a5sT+K9ddcFhekWcXBL56uLBrXR1vbac/k37FxU5Wz
5XSOZfRPw7Lr0upP+3OmqXvJWKzvH/FxX828FBvmi3KEckUejAnyFwGldPDy6BqafqXAKbYrk3lx
5ufbRbzVepTRVsJlXZ9Z5M6l5WJ9cFkavKQG0HhLf7GL0+JfjEp5V0SAjN8IoJQISZPbMyaiOBh8
Kn0Wq1eSN/7bmmpZ0Whol8sDQJvC5Iu1leO6Nfz2+9SJjMrP1V3UI6T9F9JFDeXqZP5zpI1u+s6S
Z2MqGpe+W5owbPStJtfXKbmcEcfaaqNR1HsU2YZuWo/Vid047Bq25JfJTluRMEJ5yvq1PA7VyPu3
6LOdooq+PWr6OHNYX/EfXnoTNuD+S4ATrb9QzMYL4WCvM4Z0cpRyh9oovX3F0HVknZN1sQlkqyGo
5UorGoqSPA/BZikrjjJ5HsRSsxDJqOn5CJ1/pofQlK9MmC+KmdsfWNLdb9BfNjEc9n5LGlt8S+KB
tsMhjRT9i/inSg4AcpyAdtMNq3GwM3g0rOXgzriZb8/vYBYw91iBU5DxjvCBKhk2AqQNLy0o6oA6
YfADhi+EVaYiKQubev4LaAuk5BhZDHxM6cpNNOd7gVl+57oFd6Z8vYkj42TLWg+Nv5YcxVvaiqcF
oa+m45J6q3oUVRiXLqgo2PLShlAkKHxjrzWQhi7zyQ3dLZQJxeegxrFaPfz6RS8TxPB2DdT8d8kr
kni00tpPGmcI/aQgMZxkMBBsOQDxb9FZqWCynKvjZvrioTDoH9kOD6862ynn7HTT/nHnf05sCBkt
v2DOI8QRcOs9MfehURpkgnMIo8+ucRSs15LRcUucjcLDhW2XDe+/YalGpU/XZ8dS68+TxPSFGK01
6LoSLPh/2QFt2qwu9EI3Vfy1OJuLbkv1jO2FoL9SrKQgiQ7Ay4tLnb9lAKB3WqPYJSU4JlPCzX2k
Z7C/RYKCe7iUX64PEm2/uSFovybuXfH7vmaNXU8LqxT763PT41O4jT20WkVmje2EeOADaavwQ4sg
yehTbnj16PtsetVygJkCVhusuRbqZ5rUdfNJomaUUwLeky2t41LFwYWz5aePVPzjJGIJkBQ8IfNe
dRZ/RLtuHJumkdSmNuzhvQbbYcO7GXPJK+uJBm16LsK3P059ChZpPc/ILUOBN40Z1XX98BgjG6pj
uMrLCQge9SypRK7AbiJgQZ3XbcDgrujgeBbqI5Ky+ZSvqioNRYB5Aq+iwLN+e6GCGCmQ4VqjlwpJ
S0f/JLtEhkMJvwVEesN6VU6UKEjaknT9HfcrxJ9JmIhsBHjw9HflQWTHFDF+mMp0g5bi83Sj8cpO
Fx0sOmxe1z9OK28BnIDVhTdzMw4yefuYyCV3Hc7QbvMDBj8ihRoxfcaKl6ki5J/BxFpFhHdFocJ6
jkRq7bNIglKqCfPKTgZlIVFJdPnIwYpcZf+ErV//mckrbW5fz8iiPgNN3QICw6xyFYR8gnNcR33M
HW3Xy9RxWVlsdPgNycFol4eWm3gh2UwBndSPw7NOB5K1yw/vkLgfMXkbA1+nyBXRU5Kqy46uZxy8
6mPRFdVImvLTD43ncPsPcBjX/8d0cCKjI9BxpYK3cfXkODp/hXFn10lcIuKyCwGl8+cMQvd78hFh
pE5fCC9xolEltz6aMr+AKHehcmzQEERZEechfUr/aGBVnFEcaUgYJEDtClfTf7uENxd01EOkHSsx
iIhRCTgJl5aw98lwxYI4KfAEjFQklFppvVQpUOSbqP0wapr6+0LFy5SVYNsYE00K8Ts3H+x8LTos
aytV5HiDsjuGbKk3zJl9baBZ/4HTQrxGig==
`protect end_protected
