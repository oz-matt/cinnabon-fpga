��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o#�\ �-y�U��`�/�v��G!O������)z��E�J)�ĲK�B�j��=�M:�ۙ��X�4$jÓ�K�Vƍ�P�׿_a�fC�ć�E�9�Q�����+�v�k��y��P: B� 0�@�n**�{��Gе�g��	��2PZ쁬�~���g��0q��"���x^;�o�#S���C'n���$��69�Vo�؍z�b���y�|Ҽ��;$�m�/3-��b����[׈O�����_������Wh�F���J�Y�O�W���Xw/.�j��5��sUН>��y�Y�?������?l	�vB;��L����Hj.�M�!��0<#1��)�P�eT}4���B/�N|�t��qz��*������t�����z�^I���$E��ǡ|����]��;M"Fcy4�&�3���5�����)�f �`����/�k����������A&���`(0�I!�PXⲛ��]�G[oP.��7������O}ۨ������[7�x!~ n�@���=Eꍽ�T<Cn�O�����8��Z�a\�Vs���9��A!
�g�G�e �#XwM�J��xz����U̹0��B^��S��򽭑W�)�U)kP�㍆��R��vU5�5�e!�v�CS�BD#����f����|v~�P2W.m��G���	*����N~��^"j�X؏6_v�,y��£�m���������Ƣ�-������=&�C-/�k=K������8�>Ɋ�F��e�A܅[����'u�;�1�xͤ< Xv ȃkì���NG0:N9�!w�4��G�"S�Y'r
W�
\>�|��ˮ��|�k�Al0'�v�IRu�
�t�i���H4���l������e�c�'�s�0�y)��!�a���p�A����ی&�#ן8B��%B�ݷ�庙)0���Cq/¿'@4\`�f�h+���`슎���?iϢ0���� ��<j�X���3�5�D=�:���$�V<Go�r��X&YZ{U�fG��mGVd��[�̞��>hv�B�?�.��E�黬��M/�x��y2�[���A!�7��;�49Mbҷc���r��o�§!Ь�To��0&�q���|f���+Z�� ��� �,Ӕ0��
2>��>i8[�X���Y.�.���6��."�� Ǉ�!|���v��Y�栃�]O�
��Dh}r�L�M_��8���U!�e�{���h�e�Q��V-��3ܿ�Ao��7���HB+x������������a �y��$�F��C6s�z�E��%�m� Vrߡ�_42�����ñx|T:��3���V��0hTf�ԭ���Շ�:��,� �W�����@�<��'9���ǂ:/xt\�A�}�J=Q����N���[��S�ME#M�Oz�s��[	�?r�)�/��bpi�J��E�,����"�I��Q
j���H���Nr+�79�j!���)�/��7�"��lm6�ί��<�|�)���4e�fu^�{���b�֧�
�y_�|��^��%Ӡ}5�d�\��g .�j�`a�w�h��)��u���%uZ��%c�V-:P��1�)z�48�/>e�>y�����N
�,���yנ��������8O�Z�-�3 Y���f!�yŨ��S���c%"n=�O�!E�+�i֓x���?�x�|�N��G *�Jy��ҟ��g�G�(���n��]�6[^
f%
V�I��ɹ�G�,=`f���l�T:@���?Әp��
Uy����bc?��`g�&<�?�)	O���p�ڒd����ؚ:n��5����Ǘ�U�i���s���:���HW��8�;],� �����qS<Գx�s�+
������cǊC;�8�9��Ntp7)<�i��5B\U&���+���9ΚT�����Vm�ZU�g��K�$A�d�t�L�N-�w���)Cw�U��(�25���y#B����(I��u��l��[)_V{0A�"�]��������c�Z�c4�rZ�'t���dad��D(���v@ף!h,^oӲ��b,��SA�����K��j��"�3H�,oe��������n�}-nV���a����n�T�$6�T~��H��[�V<��F��B�I.l�*I���*d�DZT�U�@�ݧ����$��atK�b+���Q������R9�b��	�!f�uW���S�3��*9��H�S�%h0f�T�S[h�L����Z5Kl0��ԉ��<�6�Q�8
-���Ye[�[m��?�8�vօ�ϿY?=�M2���C�2��B 3�CqYX���S��:F[�;�O�f���p������+&��
�W>��,��1�|�$l��6����0�Ɩ.3�ڈ;�h���]�l�Y�*r-�'��99�=�꽟S՜Fq����T���Y� =V��Ӕ�e���w����ͽr�|�
q��Awg�9E��jn����0?=�g+!FWu�H��XF�9V{%@>i�5;)��+��T�a��w����C��5�r#ô*��:E�`��[k�u|�@�Z��o�qc��A2?aUZ<d��D-�T#^k��"�I�x9G�SV��ڇ�4Dv`�g�[�<�w���pc�B�~���gs��5��R�$�yO��{��u����"T1���j�5�B���L+'i�  :&�0C
�>���*��� ����!������Wع4ސ�|�Rj�$� �`h��LŒ��o�t�'�a��8��=Ą#��`�'�w,.3�"5����Y*�������i�	����$/;���^��u,qE�q��>їZ�M#!i]��+P��`i�QOA�H�/��gu\��5�j�yg�H@�-�Q/(�䁄�7���S�~ �������67Z�L��T���I��Ȍ�.;L,G�mGj�*���_�b��ZrΉa�n��g&�ޛS
{bN�l)4��N�O�*�����u��aR��p��6�l��`�0<�G��
�:�^�E5�Z��l�&�aֆЊ�([>ܿ�N�C�O��D����*���89z��
_�3T�{���Zq�j�Aa��h�T�s��N2�J(��P[R:�R7BP7QC5\%�j��X�O��i�=�ŦH��|-�r�nx��>��l����!��Ҏ�jT�>Sɦ��(%��ε���8�FA5m^�C�
bŹBxm�#a*p�e�M�|��=��[�8��������f���^q'�G�J��3��3�丬��H�Bd9J�k�� ���,Ov�Y�h��Cl�p��2���*������Up�#`�)����?����7�7���n�e̗�������d��H%�%aK��3�ꄥ9����Pf �Q"����^�d\Ə����:���(H�4e�^�@=d1�\���Dr�L�ڕ=�z=�CH΅)O.6R��5[/�r��-�sH��<�4�J��'��m^�
�}������˚"H��:��<�%�;P�Ѵ}<F�q<���ZBu��bk
��<����U=�'������b�������R������'�w�Ư��9bk(��u��e�X��>?�a�t7�!��G�?y���3�{��>FN��ۈ� E������C��f2h]�ՠ���'>&��:����Ϙ��~ez�Mu7&�@��KA�� �տ.
I0~�-BƢ�p���A�VR�,�i��~/D�j����R�)�P���=c�L����45�z��k�9;��Ei�`ې��U8dז�5���#O���}E�!�zDy��,!v��:/W~%�G-u*
�U�p�CT1y~���vY,X��^I���8�]94mX��b��H>B0���r����3�qȥ�&E1t�2GV��PJp���ü{�ݑ��TY�1(c�Ey<"�sZMDlK8汽/E�?·�����=�Tpv�EkR�J2$#�R�yЉcvj�6~%9Ǜ��U�WIçz��d�3�#�;�J���V�p�nJ��)䲠��dI�|��ʳ.(i9E!��3����H��4��ȞNeX����t �L��gExVI��*pP�\-{��@X�uC�Bp$����D� ����d��af`����Ӌ��B�D�iϨ �戵����ǻ.�x�O��W����΀fs�檃&��h f��2�g�+�T�{��f��h�{W�=S����x�}��h�u���h�+�F��O2y��=L�Ἄ��tx��V�%x�J�8���	�N��Y>�.t��ya�5]�ޒ����.R�|��>]�tO��;�cRP�am�5�����Z?���hA-��^�qO����:������DY�W�fE�B��,7�R/+��g�1Q�w/��#}�X���=v���'�_CzV_��"7K|wڭ@��J+vM�|��q�}�x��C�~'EsF��p�n/�,/Q�S��XJLt�"Lk�%�z�0�+-�4u)	*R����So��i��0�F��&<#X���S;�`��kZ�)8H<���y`7ο_f�� Q��ǟ]qB�����-_�||���6iR)U�)5��rʮ'��<���^ѩ��%���߫��<��M�9�j[dp�_I	��N}D�!^�hFT�W����g4�l}����(��	��O˻^�V��뫵p۽�z�b����@.1=�Pn�w�)���Ϩ�4�v߬(�Ӿ�@� ʸ�翈RFmk�x�"L��S�Sr�ET�r�q+ׅ�W,�b�gɥ}��H��]�6q�#ٻR5��k,���;���n��$:�t]��&!��E��;&��� >�m��;m3��ӧ� �R_�k+V.&�՛rp�0	B��u�6�%���p��f���g79�#���$��'SK)f�+��H���^��h�9��`�sya��MT�j�|�C �;�u9�i[Lp�w7�vE�O4@aϖ� #�ci����1�i�'Ʃ�-[�fovon������N��_���*�HTL^����LW�rà�X�^9�0['9I�n�O��TV�u���Y2�{7���G�4��p�p�`)�k'r>�`<�{uw1�S%�c k\�V(��ct���m�����k���t����?����c�\*f+1���j���3�ςf���a��NT�����tӴq%�Z�.ď�Ly~j�k'|��Y���#"t��������L�f*5�n\l\�a��y�)"'��hT�mW�ε;�;dA��뉑d����/�R�&U_�[�5q(?�0��`N��A���9� �������̩-���ר���%s{0����I\�2m�<q�o�j0��� Ձ��xr��Tʚξ��Ւ�֘���m��ؐ���N�Hїv�l(ɞt �od�Ѩr����]�{z�-���0�_OƩ�.5��O{v｛�b��㷏�?��=4"�fM�'�;7�ǵ��|ns����sr����k���v��(4N� ����ڬ�q
!�*�V�u0�#��!�l��	G�e�ͅ��i��N��c����`��.�+�W��7в�V�I�\�ߩ.����G���� �Y][�n�����pjD�z� ��i�^�g1 ��}��m�G�1�{�ڣ�[�,�hK�ǒ
0J�L*������!ɞ�_� �K"ﭏ��Wjy���}c�%���Fg����J�j� ���DfTҊ�����
#�C-��w�I��N��=��#�L���5ϗfϲ���6��2}w��W���
#~h�xR��5U�lR8%(���� )1b�{��f#|�fc��G��k��`���cy���I��M�����-�q:�Z�����gO�����4����2�u\JVZ�رę�	�8Od�&�$S��d�8G>-,2�ڐ��N��Bb��<�4�4˽Myk�� �5b��ǂ���i="?�M`QK���H���U�*��-�bi���J!����K�2�J�"6���As�U�O�ޜ@j�MVSb��kkڻ��%��,����Ld��M^�o9Aq|�g�Y��'�3-�i�!6�����g�u���{��4WJ�Tmt�j��ݬ�s/(�+-G�s���0pegV��є����ÔQ�I���w���Ep�p!�L��	}.-�G-����N� ����:E�_�~�c�=������]��մX�K4o!�k-����:�7�0��]�7�U�r��+�t=('�2]��2q�M�'�e<�H[J����%è��}����5�^Ut�u�}x��ONײ�Yv���\X� y���Iz"Vn�-��+�]��8r^܈/Wf
Tv�pJ�c���VfcFG��у�ˁ��^��x�5n�x �J������^�թu����c9�,čEڭ�E�������D�X �]a����h<������f��k;��)� �N&6߿���U1��|�;�%'f����`җ�^��aAh�D����֬Y�G�Ax6A8����?��+�K�A��E�vL��'��K�>FT�"m�e��r���k[z�Y��@�_��3_�t La����EעH�ˏ
̛+)V����X����!&3�s�&�z����J��U9���:�+]��p2���*�4fr0R��.M��Kĭ��e���a��#e�O������X����E�Z�i�7aڇ��q;�Ƴ�C�Y�o�����\%i_�]x1�Ϻ��.��tB�*�:\=F�3rC��fe+�	��)��1*�y�2{��|�g��`�dȂ�x.�O߷Ǭ��.�l�
Ġ�+2����h���4�d�O�`�G���x&���"+9D��gږ!���2*@I�bI�=.{/AVHò�$���;H�d�Fy�*�i���Sk�l'��b5�����ۥ���]b.?�zl�hW���u,V~ʍ"�su����Sˑ�E1%��dNK��~�[�?�m2���}}�|9��8>��+�Vѭ'�"����C��l�O�*��Y:n��Ѕ�Ngq萡
A�g��%����;s�+E )S�l�S&�A𒽫l�|Z`������2}5�N.�ܕ��%p����;�>�s����QN05;x tu͑���!y<Nx�11-�B�Y��4T�/2���&�q��7�[B_	�:�cu��n�O�T�$I��\�B�P�VU���F�̓�j��Ӌ��7��$����0����L�e�Rc{\��R��nY�8��c&�������@���պ��Ē��6�qMU/��A�4~٩3���S�N\��~�f�|�yc&ǻ�� �8��n�ye6`'��?l�T�n�����ő
4�����질9nɖ�Om����P��kGq�>�Ǒ��U�rB='�q�j�3"��>����t&v����r-^0�⒣-�D�yH���AD���#��$���d�D3����!s���A�W��tȧ��x�g��c#�rN<��[?�N��I��k����<����h�0�c�	�u#f��{�@�}9P�=����|\;u+/y�ۏ�$���C���w�3�4u����~"��h�������ڥ6��Sټ�m`⟭y,�� ��3#��Q`6�Y`�Q�9���v��������*��O�4X�	��OYB`����4���m��?.����V�WX�L�xL'>�[��� ��e��o�!�=1t:�)�K���΢t��y��R��y]fY�)��q"p�W�U3n�7���`A4<$�j�G����{��(�j�J��Y�RrӺ7[��V&̜�3��~�nW�[���W��	5�S�<��[ZH�!�徣����`R����� I�{!-��h�=�)o��9踊�{s��W���7O���������:��ai�5KqglNFV	�PJ.;Z:4�M���0���7�i:��t�y�kи{�G_S��)��`U��(���?�&�5 ��&�-�1$��*sajA��>Ь;
��O��S�������T~	��>�n���
�8�X���  ��/�������_��X���\�����Gc�H:&�i��
z�B�)~{a�ʺ�
����{RI�M<?����%NW��-+ 6���-*1˪�_eŨ����k2��laJ�A�[zοɓ�� ���V�(j&(�JОH7�%�b��)�.6l���2ݭ�vz�W1 ������ϯ��69�Np�f*�|����Dxd�>V#�v�e�S���E��B[*�1E�.�|Ukw*�����R.4�cZˋk��3��#�;+�����Iu�,��p�������L�u���˸͇�r�J`!]~!��?~�tO��+�S��US����J��%����X�"�ԯ�G�y���R?4J�w�mУ��Bly3g֮g�3��U[�h�I�jr,�R+�_M�#W�Z��k��}Y�}g����������Rm;�Cm�f�s�L�5�@�ؗ��tW��i�#�n�>���1�N��Aƾ�X�{Sm����4�w����	?��\A��n���*}�/��Խ_h�^�"���X[�f`�[�nĈ����c{��qF'�h���v�;�E�����|�À��Lk��g;KD������bl{3o����u�PN�{zd����4n�jt1���N
Q쯙δkM����VJ�c�����z7�L$U;ky_�s��0�湕2���/��1��v@~0'��������>�{�z-,bA�L�#��Q��?���cu�����0QZ�p�-85^��>�,z	�!�LƮ�M�=���mz6$P:{��U�)v�e�>�ܮ
0�(�ߺɽ�@�Y���D��e��YE�u+�A��r���'�) ���ྼ��F�3!%ةP�����glď� �J�\�Q�z�rO�$�)P��z)'�i��e��j�͉>Nu��G��m�����8�*Y�}-��/@���[�=.b}��\� DF���v�5����x��'����g}x/��Oy�Z���к�Ε�i4#��,J�(��,!����r�r�b�Y1A�x�1O�:i+�8\m�.�� �E��"M�c4���8�L�IaÄv��ְ�b}���?�ݘ������	^@�w�OH�6]�&�p���/U@�ZZ���9�U����T� *s(g1m7��X�\y�Q�J��5�-�9�`���F�x
�� ;yK2����s��+�m�
���:��Wڤ'�m�4�	n)��i���E�əa�B���n쵍p	G��Xˆ(����+��X�WbC���d��*���lY!���&r){q�O�7��X.�Yϙ[�=F��)n0��{IB�_�0����*��̰q�62��0=��<Q�饺
�K`�R�N��c�$=Ep��1��\�Ʒ�����s�������2��}� `b�E�G7��)K��:����c��n]/�jf��ݾ���o5�#���rZ�%�ŲȒ����6�Q����F��]|C)�����ц7�r��_\�)\G�R��*V�u���郵.��뒩�|Ql57&��u{'�<�Ѥ���4[�ɸ9��Y�ec`Uo�ݳi��Y�w����)���rj��_�)�
�avU< �Ep��$�V��cQd�̚���~����ir�����N���*lD=ELFc�2����dQ	T��~�k#$:���F|�y�ɪ�!%S�徝Q�H����`�%tG��Cl���gA�ܮ:Eq�n0�.ǋ+�3�Z7Z2�����U��n�C�~s����9A�L�D�����z�����1��U�j�}At�>�Q��^D�C���@	�ʾY��g���Ê��T�H6�2&�9��dk�5�l��dO{�������WT�*B���D�JBg�6m�%=_��%�M�^2ծk�ݓ�>��+�ײ/XQH6^������Ѵ���t��,��ݿ�F%�/];H��P��ɂ���h��4T�	����3����wS�F���o�'���w�oCǙEH���(��qz\Qe#�&S{����aW��j
���K��M�:��4�{j9#����m�V�ӦY��~pI��ݞ��x�!�\f?�m�5�ň��~�=�"Zh�5Q�<;&�Y�,�姕G��t���Z�V(`��~��RM����W.�s|��l��Vmx�~o���fe	�t��Q0��vx�X��I���3�o��1��)��5&�ri�k�j����X
0`�F�{��/Xg��6v�����t�w�dP�@a�� c�ÍY鍆�^�j5kW��B��;vϋ�E)�?�q�)�C��y�hf�S������9�rظg�6�FB�?�s�9;	Rv¨�����˸��$UZ5�V9���|�-���T�f%}ꥴ�W�ꉐN�S�b��-�KTF��x���k�0㓢Qx�[��Ih��V��&��q ��~��a��_pk�;ϩ��Z��8L�k�[s8ą��(�����$O��+K�%�Rny�R#�z{��Q�M�G	� Kaڀ�y�Y���?=�����`�m1��s�k�e�b���s���9���{���\��"KAM3�Q����Xu�d
����+՜�=�
�v��}2)��˲����;��~F�?������)�����Q��i" �x?o�	�-����Iw{���x5��|��(&B2B=�q�0k
���{&�eS�RO/,5)2�)=GҔL��z;]�"�܄$@�,\���=a(/G�;G_(��PO��o֜���4%c=&	}�H�4��g+̄�������I\,���;�k:������i3j5}4mTU|���|.���d#Dey(�5a<��+�bH���3�D����F�J�9��ϭGZnDXM�p���P��O')䏊�`!R$�DO�K�X���Ҥ���?��[���g�"���{�	��k�H������$��G%+���:�0�YXbvG��iN��Rd~#
�.M�ݖ�KH�Z̀���gI�jr]�.�?�de.Q�aM)�kI����Wc6G����� o����1c�Qn[�m��V�D`�d�=���Y��>.����}��ҕ�Sh�k�&J� �O�1��Ju�U�Fu��<��d��Ğ�?I��D�^�{6;So'�n!�;3/�}�jc�8+�q�4�� �:�@��	�Q!���2��%}�Ss��Gx����Z�H4֥����B���GRb�uj�uu{�b�|����@K��K�"�@q�m9���� �-�"#.��F�2D�B�ej&�z�1����I��Eݮ�@kj�TX^b��q�����x�cBD,�HB�*Y�2v��5v(,�@їz�$T<��۩��2��]t������'J;:�w��f ����rŭ3 �B%� �ʨH:�tiX]&e���B���`��K+E���ħ�߰VRE	i,�y�m�EK��M�t7i��vI��Qp���c#D�׌4��?sF ��^������Lp3��p�WH��%J���=7`�!���TP�n��C-l���Q��<@���*X�f B���n�PG��Pi��3�`Y\T��{��D��@J�G�_;>T�������}�f7�赅��N�sM�{������l%��Mꕇ��*S�E�h;�g�$�y}NSy��`�-�Azh�i77��쓹��]�*������[�Fk�����+� Q��253n7`A��\g�/A��[��
������Y���Ϝ���1�/!�_6gV:��R�������'���@ɚ�]WM/W��Ce�X Z���qz���=#pa+6}���N���?�|#\|�F!p�ԃJ�;s������=d����)�!�~ݐ��A�G�N�F/Y�^"��:��F�%�\� %�xޙ����0(.�g��]��K%	#�c�]��m&�\�Y�u�ܸ�������-U��@jg�g�����E͙�p�/�E��c�k��$�c�"��������<������i5]�6\���i��-�g!�@v�=��Y���>�	.�����1�ċ-�����BFc%�,�C���W��O�c�˾�q>-��e�O��Jq�?3K�;�>)�n�%����Y��JI4?�Xg��%�Y�� �#n��v8�Jm�M�/�0��G�v��>� �d��z�Eqb{5�G3-��$)�Y,C�lG�0g9��,b�Α��s3$����c�hL�)��� �^{zT�������GԬ���T?M��^� �>!I\�q/�!���锼@�Ԍ�iq���Μ'Tk��w�3��!�Fɔ��0t�;A,?݆s�#of�?O�v�c�%�a)d8LdaA3�,~[�,���V�%�^Tӟ$k]�C��b̘�8W���r���D�����%� ��O�Ȧ��h�ӑ����&���y&2�i~P��hk^�坴��_>�hG�h�����wH�ה%<��ۋ�ۉ���7��	����26���xT���A���X��b�ʤ�6W�qM����?��Vx�/��PX�����������W���ژH_����.�M�� �&HJ/�F�6`�&�����K��!����LW��:����ȕN�j7�O.i�0�2F�ߎ��+�q��M˹��r ��ee[�ܕ�x���v����iE7���TO�8����H�����6P��S�\�8ԏW$�#h�VC�M��>YAb�h��6f��of^�By��4�H$y޽�QvI�S|��0�����5��_�R#l����H���T�L�f֩v�T��8������ \��"ڲ|�4�ƽ����[���y�8�4������H������9z����Fd	O4�X���:;�u/^Wuu��r�J*Z��fеu�yCe�7b����\�����V�L?{:�f�ZOH,��^̔k_�y��?5�]�T�� �(4\�۶��(}��!�|T6��N� ��̏���;N�Z���"�D��r�^�hڠ��.��R��O#�|�36��f�j^�/�Z�AI@�ƯI�#��'������"����,�9��)���$�{�Z��g U�\�}gt�ң�:�F��w�Ai0)H��y��@/�؋�~l�Jr�tt9��G��x��YW}��M�Vh�_)�Z@� .d�~���� )�]q���f>$�P�#�V�<F�ѻ�]*wϸP!P81ad��XO{���R�8�į��E�_������Q���R6Z�7#��Uh��
��x5�Tyd�
�-j�mQ%JU&n|�=��u�n��Ƀ���%y��y��n�!���/��O���?�z�͒��x�tR�y�P�wk�O��9�nKmGk�!�K���������|�R��������cyn)C�NM�.'zQ{��8Kw����ak�/.�]��l�g\�b�7n6�W0�H������`Y�b�39������S�_�[3�ؗΓ�/./��i:�R'�W����>iPK���+:,��Ŕ�5M�5x�F�+_H~�n��͐��݃�Eq� 9	j`�W�ABo�ZP��ޓjmN_7�(ȻJ��rgQ [9 �t- ���(�����B�#vÈf�M�I���<t}r���7kx���gH��Xx�M�GZ.�ae��*�d�峾B�+&�������I�cC�]��SC|�����ؼ�G8<��L�JI����{�)�gCXӬM/��2��x�
J�M��n�Ѿ�.�E<��1�¨2�q֟��V��*���U�5���m���Y*wl����p"�u�H��ue�֖���w�����QJ/������օ���،��?��%�����y��pmO�fjE�5c}��x��&$Jp�nյ|&ܫD���ʔG�|�K�fT�k����U��C�t�:Z�B'�#hIe�N�0،yfO
c``^�t׽��O�L��4�)�FA
�5&�IG��#�b�PUx��;y��_�PN�dx���^U]- v���J?�ϭV�(�js��������a}(��ғCc_�f(sP=�.pݚT;c]�?E�bp��P���<�����e,�9k� ��T��-V�9�ŀ2��M�=�f&#ޒ�ib�� �,2-��������n���RO.�X�	�%e`;��S��>vۥ�\��)��ሟ�O�Y\w��Y�ڿXo j^���}�ͣ���I~�~�c��}y�!��ͽe�Z���!�e*u^8�����R��Z`��G�
$F�����7��kE��ahʌ׍㕹�* 2TY.�݈�^��p�s�B`kj�U9!4��3�É�������5����B���5+��J�dQ{�Z�O'0��A���"��hp����sa����b�=du������at�g���b6���:�`,WW5�:�[ݑ-&Fd��?�a��*gv���R�����1F,0���[��]NF��l>���@�p���T٪�����������-�ga�\n�sBb���bn�߷f$6!9Nn+��O�L��x�x�Yy��;���C�q��>Q&�t���k��WG�g����|)D�I5��w�����[X'b���P V��A#l�O�*�$�t��W����L��Y�-�Wv(�����[UZ��M,�/��h=�}�����'���1,��J��<�A$�|�=���Q��f����N2��GPO�?��G�d��o@
~9�y;~�0��	�:�6yȍ9��5�.��G39k����x<f>`��3���ߎ��޳���ۭ'�wj�zu]¿lZf,�1y�R�q��В��g�Gw�ͦ���,3(�5ϋ}T���������N��,��G邔���K�G������W�(�3g6݌���P��B��{F��_�����4OQз�4�w���t.����i^1�Ӛ5����,�>X�k����)�y�)�Y�.��Y���{�01���k-�0�Dư1bx3N�S�]�s����dw4ˌ42X��Φܢ�j~���z�Er�+�N�p]��9�w�I<��l1��tS��y"JN�Fw��S�����[�/�1�6�X-7��� �-̷E8�j��>ͯ�Of�;N-�T�1��0*0���WXtމ�݉���8��Z���a~�����o `«L+3�0 Xk�Ki�}��G�Q  �'wլ.'�>��4dze<��4 �D)k���-g��y6��.3�aiei��.��;�,�ˍ��V�@�	X�tqw�<�
��X���)�-*�I��xkz��Tڇ�z��0L�G��՚�&\�7�;m�F`�}J ��o��p��#"@�qN�|
�(�`Hi%8=��[5��jml͹�����V��,4l�/#
�������)���(�F�����|�'@(���R�y��4�WƉf����xTa�n���o��3mYWm>e��Ƶn�Ժ��<��8T��4��d�&�=tJ�0(qA�e�Z�3߁%�w�Rnm����Z{W����K�6�F�,>���x{}�j�+3L��o�uB=����k[a�����O`�T�/KҾ�u|��#�z���\�\ ķ��҅��2櫔�L�ϰ�5��2� Q��F�`�<����m��X��zK$�r]��7�=�s?�E�h�.����[�>e0�����ĉ��p����E��)f7��"�mV�6rx�-.L�A�*h!C�}c��I��9�`���Պ�p�]�M(=�%@�m���0�f���3�A�I��)�O��Չ9|����|)�b����އ��8��pQ@���w�ǵ�q3��V� �_�e�3��h�f�)���	lώI�X���uB+�kÔ�U��Y�czĔ8��܄���,�#�j����+M�@����Sݩ]k��w��R�w�n9"�������"d�w�L6�����5D�2� �,v���l>��APX�L��\�3�*���ҪG+���v�9��V�����W��w�bW�cD�����ņ0V���/B7qM;�k���������kGm�$Z����3���t]W*$�>�B�o��#�`�΋����r&��-�	h+�AxW],�Rޤi���qlxM�G�� ��(8��T�  53����?	����*hf*o\LH$�1O>m�e�%��C'�p{�u�� ���x�P��,�Y��ێ��Q��W������t�*ozN�jH�f}���t(Z������1D���]�:�����8��o��H�!���g\����A�>��s.�yvb�f�U��D��}��A���P��J+J�3k�Q�Ag�����qfo:F0�ul)jq��3�NB��:Y�V��_�+��.�w4̶��T��+�{�d����:<}�5�/N���s�ǂƃ���v�U�)��*�K
�T�LQ�x=�_�u�n�;?�者|_x$겧�Pi��JC
]z "�O,��� ���w+�6+'��U���j��-�l?|
��X�fS�;�g(�$>�*����V	������5�"�=�2z�8�����z �N�9�Ĝ���!(�f�n_n!p%�LT �b�[�r����	�`7|9j�^��H�/0#/�+3II�Jo�*�,@31�t�@���{9U;x� &R��?݈�s��"B����.��Ȥ��YĞB5��r?�sK%�$$J,B֫�="����b����~k
T�N��rhaD�Ϊ\��8ն�Y	&2<����$ �p�26{?�i�� �H��GdÚh��Bj"���Jqt?�8��m�2L�L⎹��\iT1"���-&���C����K�Rh�a\�x+���4!���U��Fɀ�:Z�2���9S.�uv=F
�^�Y�s�2P��DT��ɀ�
�j>�ȉ�i�ms�c|�f_�*�6#�*1盼��z���9�!8vUd�aO$���9&ȏ^���u!�R�4�NC��KB"����HF��.��/�!�k{���4��[&���eE�䬄�Ks*��	��j���GG.m#(k@|îU�f(����%ߢ+����_,�������*�M���U�9z| B�տ����l�rz�[CV8_7nz�w�q�x��V�$��\�~�
eM)�n�&���
��*3��7_�I�%1� �X��^�?��Y�����S&��YS`��{�.�$�%�e�]�g�^=�#�d��a+�1�_!�v�R1Fn�;~��T�ѻ�g�zܭ�
��QR���WZo@6s�ɟ�4��m|��M����և_���/�e�"�5<�%�I.��i ���2�C<$� ~�%�������v�5i����RL��~�i7@nw��+f��_*!TS`L�����0�RZ��A~ih���r|�LQy�lS�ʍ�e)���^8�����62^8���#]@��C�ڤ�YN��H�!5SVr(�w�y}�_�=���Ƕ3�3����:s�~�eJ'8.��A�����kũr$���*���a��,~��p�qKw�'ɲϵb��`�����>R���Pg/�ײVa�?�S p �������a'QH�Y� {����_8i�f�*�yJ�r�%�>��(B;I�[�E�%¡Qq�jIK���X�r^Y��=>	��~�HC���E��|B��xyl}�8#��p���D\W�����ӽI�9�V�
)��x �����T�fH ���ʡ�f��ێJV�����
B �e;�\^ځ�m˥5�̞Ce7��0K�jB�W��2� ����L�8�&��O��A���eF�/P#;F�gd��G��[nTV��Ë�k0��ׂ+�u8�l)���D���8�d��S�:����| d�%6�_��i(�n_<�>� �M� 	���o)�+��ohD�A�gLVnL����I���[��Q bk�xC&i�����j!��D sƼ9s��G��q�.#9Qw9��ܒ��A�d[sD�Y�����BPO;��@g�2���2ooW������N�H�SAG�t�nS9�*C�� ���b�٫F�Q��N4��Ab�c�L���Ozb����k|KEn��\�e���xz�n�OP��_�).3r�<<y,�7=B&�`ZK#���L-d0ml%���$00�2u~pW ����5���z�|��v�_����z�R��]&�o��1P�������E��I�!�����Gr�E''�:�*��x�tr��G�s~5�ҊL�7N�++��f�Һi��V-0��<�c�$3��)�zKW�"W��be��Ƭ}=*Ad�,o�� ~��F)���`����
����Z�}�ۭR�:@�+җ9fp�,Ü�� �z���y="�"�{���uH@i~����d9���'�pJX'3@_�*/[�]p� H@�yBU_-���!w��I_:KM;nw�1���/H5���ϩh���-��w�U�k82ݫZ����ʋ]�� �qi�~l`?��5� ���ʉ﨎��{��`���Iń�ya%M���Bۮ�������z8����05S~M��'>�?��.*B�)�'�[���-C�oP�`�[%)�h�B�&���S'M?�5��+׫�\'����PY��=�}[!�Q�+�֜�h�v��t:���#�����$/�%��M�t��:�� ���8s5j�U1���������uނ�ߩ�ݔc@s߳6L|hg?L�
����Pڧ���|����;jg:�:���Թ=�#��x"E�?��8�zK\n�;o�Vn��٬�@'��M�V���El��� nwt�ґe�:R�{�&�B�j���y\йזj*'�����Vb���sQ'�j)��X�$��Uԥf�8wK�kJ�>H�-7����fpS
nlz�;q����:���[-(-�������!C�,	��ա��'��������l�b������\�*8Z׺�@�ӹF��h�ּ�!c>?V�$<a6��=��qG�EX�C6���C�Z*:!�I��t�pBE2�IQ��O�eZpt#n�wXv���>��匲A�߿����9��i^j�6�~븞��Ǎ�*�8��j�|��Iլ��������W�"BE��]?M�хc�O��8���R���R<%� ���* �\2����$O��q�����e0Df��F��=���8;O�JXN�ES.ѽ7xXgwx������,�W�EFAo|�`�y(��������g�_���&9g�-�i�v�3agC����O��y�ZObED����U�-�N�i�jsK=+0r��ǭ�kھ�Lh���y�ο�HD-�@V<ɬe�n�����ώ��<����U�T��������1Gȹ�〰��E�n4�j�^B�.[Kt��|��p��@̸j-|�<(�����3�p� e��l�34�Fz5�6�e��b|�^j���a�l�X���#��|�+#�+��4��y�4�b34�B��2� c2%�U_V���&��tT��Q���s���WB�H�2�ix��C]~��	�ù�g;���|��p>�r��� �F��E��.�	�Ӑ��V���l�\p��LN	��$��rq���7ԇي��`�9@j1�V
܏]w�x�5��Rb��;������Q\̓��H#+�3��b�:B����Q���7�_�`�P3d�8��M���9�i[�n��M��όN��]߹��P�����4b&�χ�L�������?z��d���;�&U�f������_�2]=��Lb�^�&6����V�����4@���ޡ�l���dZ���Qȸ��oq�{r^I{׬�3w�<�Va��ݔ����>��n���|P���
��(�CM`A��Z������$�W�a�OXx�q9��ۆ�!�Ugi�?�dVM˶��	w�R
*3	6�Id�t[�3q�$��m��<���E�����Ƚ��b�KD����W��i�(�D�O�N���4�>�kW/��}v��4�T��h��FcR߂�D�,�CH&��"����5���W��p!��	H�eS�a*�]��L��'+�kΕ�ZD�S����;A��#<�V�
d�z5Ð��D��r�����!v�OӖ��*B�80�~��wڦ��NmS6UQ7�e�����F!f.�AJpF��l!g bT6�^Ռ����eui�q��b
�Ld����'���k{��C��~�x�)���]>�Z���
}�e��EmO�<сYE	�fӲ�R�qEbމ����
E�0���f
�E����3bׂl��$����s�9/a�!�ؽJ�x�*��ʹGV�Č4$������e�4����;�3�h�����-��t�h����R��{��v#���ϱJ�^�%�N�h�9�&�+uq0`�i��.aձ��.I�c>~�h�XO}���JX�aG�qezfv���G��?P���u/	8�'J4�����5��{=��ĺ�,�#�~��}�ץ,�U��t��b��� f��[��f�:��sܿ��6O�*�OLa��î}�T����-�?7�3N�K�Cx�iU��\�%\b��fq��s!?�}w�B��&tu]�1�3��h��_(�2XO��%��il��?J�%�����n�v'i��͠�3��_����SX�m%�IG���
G[�O�=�����k��Cc��d�q���KAp K�Ջ-��� �Ɲ�ڟ� �
�=��[E�/���Wb�/qpb���cJѧ�N��`u�_�
1E�j??�}��%��]�_����C�ݭ����ݽZ�8�GO��Y��s�]x�/{^�F��[ԭj� FD����1�z��NKsB�J\��9�����@V��)`�4٭T�d*ĩ�[�f�'����ppŷ�WD@{�����N��o�6Lz�>#}�p#��d��`��fZ�2.Q" �����j3�����#�8zD;
�\MC������5�ݭ�?G�msfa�\��Ú7�z2&9-k9�蓍�UC�z�{���%�ꯨ��_��C@����qd����]s0a��	9�� ��QL&t���Ԣ�
������j;��(�4�G�oi�=F�'��[J��~�[�ڣ ���E�|����28�m&���O�H���ܠx�7>�Y�
}��g��x�S!h�����8�������0{�k<
�fm�v�\�+ԧŜA%�����y�5Õ��m �ˀ������/����f$ow�E�+�^�ϖ��1�P�I�ѣ�G���ӭ���&9�r���S�r5-gd �ץ:a���m�? 웈j&��� Zn��1��c�?�E�����ߥ�:�ٸ�r̕ᱹ��3�֢��@�Oc�S�����ۤݩ��H�r�A*�Uk!j𺗑� Uxl�ĕs>K��K�M#������M���J��T�3݀\1�����7B�l�.m�����[�NY