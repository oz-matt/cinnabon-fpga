��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�����)���'�LR�G��#��[,�{�̐;_�~pn���������ʏ��˨�XЊ9SF^�O��*Y}Q:[�4rP0����r#�)�(�X��"�}�x��9�e�&��=���O�X'S�	�?q�t��t����=؋�&���\��u�qQ���ed@
�l�6̈́���Sz������@X�����UO���}���v�l�+&,��I!r��"r�9�&.�6AɁ�CNS�ln�D<L���������=�/DI����ὒd9h�H���>Ox��@���dM��Ahҵ�,�b���&����&����=�����lj
t�@��?ul�n�V�)'���B៘$���FU�,G�w�j5c�_�o�F�H�- ���}���?�u�7&�h} j�
J6�b�|K`ǆ��v���zږf�V�SbZ�_9����F`�(�m%I�Ų�Z�E��:�A�gW���V��vQ�"�v���\���5zE�5����%�lc�,���G�Kf���ӛڝ��R�����Ϭ��h"�/�1O#���#�Cż��S_F-Y��������F� T�i���k�������:�Ϫ�X:6�bDg����%	�,���5�Y�b�2�7w��:����9Q��� f�������B��f��-��/�Uudk�p����VgL�cۀ����'���1�O��R��t;{�m�P0�2%N2��85�-8 ��%䳚��e�r�zŜ��"2�o��>����4����Ɓ�, �^N�j6��E0�;
�n�I:�fZ=$6��G���l���3 S��,�i�#>�b��(n��7?n$���KNi5��ͅ�^��f�T1uo�p~JΨ�z��Z&�C��x�":��_=1(�,%�v�r�[k�姮��Jsy�)v��E<c���E�ſ�|�P���]��B������6J���I>(����ЍP�HYO]�/�N9;����5�+�	LS���(�?F%��N�>F~ZatǶ���P����_��'����sy�ta��<��Q�X�s������t����x���*�8b�H}:H� �7��jZ�a���k��7�p�ßC����&0�$E�"j�t2��^�Z{�N�vm������z��g���2n�?�3<���i#�>6���r���if�&��_���#�U��u�ul6q
vb�=��@ҁ3-M�֞�?*>������x�b�Nh��՟���$�g&�9iY�T�6���Z�uu�M��.l��$��QX�o˩++ԮBՍ1izE__<{�����`�F�8��e]��qL2����QSu�H8W�`���w��Z'�1^1D;{���c�!�O9�Td�9�E��S�
V�g.�9����.G4:��'!�F�����/sS�, 5�t�3�2��¦y,m=6�2��S1�?�qI��k�]�@k�8K-�_�ON��4h�Du�OQ���;4��S��;(!�L�d�]�����B���FZ.�\���µI��8#��L`�I`Ν:�YnWF����oЉ��]�8WS�~�C���%���&jR󙘈CE\BgM9
<�v�9��w4K��4�8X2sB�
�%�b��E��‗g�6�v_��7�����ܫ[WGWk�0^�;x��?�b�Tj��f�x�9�X�`�΋�5(U�`�0Θ�����ÚZEݱ��pPowi�_��{�v���}�j:����V�]�1J��*�
h�N����6
��XD�팰��{���-@���ϗ��r���L�/���2F��ڮ�ti2��A�ծ�$&�e2�A���D���d4oRW�'�WG�����6y�)a��]&�OP0�o=�ʻ*E��+~��`��z���b=��Y��!G��[f��㳦^ގ6��))�G�\_Kj/��d�\6����r![�	R"����}&N��K�r`�[�X����-Yh%���'��a������/��Ў=��^ǈ�豼Nkލ<�!����_~���E� �V����8���`�˙�d���@�h1�R�#(u /��pc�3d�Ś
�Һ��q�m̘Ԫ�#|%L�>��R_�G��]�_��QL�X�*X���w\<��4�J�\�@S�aj�x����d���?�.w	[�iM���\A&tJ4/]�0����k��EoE���{��p�de��h�+�F�JS�H�Z�,�3-$������� �0�&lR�A�L��<��b��ڜ�މnp&]1�W��X8JWhJ�ֽ\5dT���-�ف@� ,v��S�!��u��}�^%`ܲ#Yݔ"ٲx�!�{��6=�\��)�K
uO[`�W�Q�B��O���ql� lq�gI� ;�5OЅg	^8�%c�R�(�*Zq�A�Y���
RZ��qeH�������:ͦ�~��u�۞`�|��Ҟ5=�ޘ�b��	E�b�a��/�y.	4'O&��F���9<�`��xB�,�s������6�x��`]�~E%����V�	r��e�}�7��VUi�^�ߢ�(�*dɤy�=�/E�v)�,��O8ߓ��2P�:D*O�	�:^�˯��ם9����v/���ۼ+�����'r��R\v�/ի�3������r2��4l�4�_{�n��L���RanL������~ﲗ�02�~��l=H ��@��/]�*�� %�|��j���y9�m�fa��E�p!dä)"X��	߇����1�f��ӫ�x��V#�'5������_�9^{�I�;��G�v��t��~��Q~��-_"���LK�G1d����僲�"�`�IL�ϵt��t�sY�Y��֔��������*,�ۇ���T싾�p�ώiW�"��		P뮀���mr�p�;���2e���bpl)��R.�#�M��<�j��Y����<�"�=v�h0�+֤�u~LzG����2���i�S3�q�^���$PϢ��%�e��z�ݢ>�5p|ho�?�/�*}i�++9W����T��Ψ�bY�hz8k���
ft��2�Ly���{M�H񾝑 �o<#1�(+�"2W���{(�s/>������o���Tт�,)
M�6�8Z��Rv��a���n"<�Yw��Q���N�	�+	��ڽL;��t���(b�K[�����c�QH��L��`Y�.B�K9D`��ֳ&E�,����Mů�t�E1����/94�ۃ-��8�G��V6��4�`[�V;��z� b>��b�<�_��Ѷ�V�M��$�ښ,�[��_�Èg6:ˡ��
�6���Q�5�+���;��B�0��Z�)�ѐ�|�"�^-�>��6�w�S-�@G�9�[®(�����]�Bw&�U7����Ll��)\1���Ax���tc'h7ﮥv?�~%�\>LLåu�r�!��h�|��N|1�.�p�5Wǩ=5D�5.����>v�%���)k��ӵ��	Cf-��=��/� [����k"�K�o�پ5��/֒��S�Ŧ���w\_�ƌ�OL?��H�Ǣ�tf۴�׀�Z�P��>��xv[���o*'K��:#D�:̉'��/�ח�H)|�S�q[پ�Kc�ZgC���������a�����W�L�mB�(>��PI��W 8�K��*[� %}������wx�"�����s.^�7sMj(�ye���m��f@? �CTa��9��'�Y�vٟŏ.:Ph���n'���Ҹ���O����Ȩ����s��9q�C0*.��I�6^_����0�R���J�ĳ��>�trJS��Fn�%%Tz�;j�F��Sb7���X�"��z��c��p�mߚ�;��ڏ&}'r���Pu���йu�^��G\>��`�u��<Q���,��_U#�Ǟ6/B��6-�=���{t�q�f�5�G�y���yJ�f�E`�	b�um����l��0���.�K��A��"x���i/ecY!N����ȴ�j�OZWy4C�\�Np�(S���9M���pS.��)��	��s�>h�f���UDY������[<"-#�?m��{�ayX�>����2k8�A���\���vR�#׃['s,��n"�q:�V��ob�^�S
;
��D��_�dc�l�! K Ɔ� e7w�<�JM3�{0���&�Nz9�p��۩V��K����vݿ�㋨��8Eh�.��������FG.E3�G]�'�]��qt��� �n����� ʷ~:U0S-!���/��� n�zE?5�j���*+K���W�������8گ��#���],=+s���a~����h�h�;Š�h9����,�������B�DZ$$(��w��5��C͕[I1���49�ز�qoՆ鴗�h5X9c�2Z�R�JZo+��L�)b;� N���1-p۫8��S��qo���ȶ9F��JEy�T-
n���4\�&V+�x~��6|r\bdH�H �h�i�H�����%�B�z��3��>H��9
"im�!2Pb��~���Q�(�Ъ"ĺ1� �3��q��|���CM�g=�p������B�r�mvsZ�f��~3��.�(@Y���"�;���~^R��t�V�]�D�l>W�Xp�I,�Eu0���q�ɑ��iP�VUB�M�ouR�TFR9����,f5�j���S���}e6�߆��Zx�����ys�bdjd��q	#�����{�m'F�2~������<�xF��I�-�=`}O��7ѻO#b�	D���fS�p�z��~c����\lh��Q�A�+��{�*D�ʤ/�)��-n�K��*�?9����9�K��{l�熸ϯ���k�xv<@�_s �̣��5͡,|T#�!�}�&0˞k��x�(�<:4=�Ҧ|"p4J����0EB���,�{u&n�E#��x����֤�I,�0���8E I4��BVs^7š���tp{�S�	�|�ZI��ރ�nlؓ�� 6)1ǭ�<�u��'���rU������$i]�\���7�wF��������㝩S���Na8@Sx�u$�:MO�~AS,y�gհ��6����-Ф0d?.18�l"���0�����m-�{�<Ճ��Yz��7�=!���~B�3��,��)�|��Nh}��(P[Iu릱�q�L�W.�.�dc%�o3V������՞�S����Jʣ"p(�m�mH�P��05�k���*'F��lT0m��Tk�+[>.a����t�	���IC#x=Ή���?�h��08��[�ּ���!\R&�KL��Jm�
Y%���5�\�1��T2.���Nr�.��P�
���c�0�(KT�����}[J}����%���/�5Q��S0���WP����+5�=ݍC�P��|{��K�c:i5�M�7j�[(���%,�O4%��j�N=?���O��DZ�%�I� |���(�ې/�rT�G`-���g:�&|S�J�S�*�Gᓐh{�y"��&9)�7�ѐ���Z�@�kw��$�6$^7q���̜��d�Ƶ��r({���'9N�1��?����7�Y�֞�uH��)�e��]ɕ��{�.�o�?�w2\�vel��X��oM�5e�,)���9��<PV����+��Y�2J��g�;��8��5h��Ck��>����
�yN���)�bKl%]�{��u:��?�6̤l pX��ͯ.D��M��h�� �4�d ����M\S ��KD!��lP�ݜm��h����"x�~�?#	�������T?<��'�I��'�t:Va��e�/9\)N��st���-Ѕ��������/���K�"ǎH�L���n7o�`�Y�2�Ԯ1}��tC�"P~�.]�u���2�0�q����:�O�bF)ƣ�fQPA�k�I|�u\�x���ˠ��MN���q5�R��xf�<�RK,O��+�%��b�c�n�=N��أ9�.h*�Հ���r��p�c�[bG"�����r�E*G��$Շ��qޜQ|���#�>���&Qg�XR ���ەPĚR�=����p�:�1�65V����+���A3OeO��b��l��D�J�<�s>���޲����W6�X���gL�
�m�h�vҴ��D�qQ�/r�A�#�ۊ���7l�wCpL87�9�mSx5^�EF6���M%�$i	7�<j� �jY-1�|}��g�T��\�����
ƪïd�i��&���,��LU�)~y;��3.���My�ëگ򎍙,b��Ȃ�F��y/x&�� ��&nZ|e����C�?�qT�&�˝����cX�~*8r�UmL���s���K�7�'Y�o�I)�[ۧ��9�c?"��z�����^����Ă�õ��J��f��[4�m	�� �6 �N�d�x�����d1����a�rs�Ғ���K��K�J�w�D��b�+�2$�� Z�zp�a�?��dD�%�3`>s�E��^�L��^�I�\E�{�{�6ZDP0P���O�ݸ��-O���Pq�em3��\�p/��}h��vޜkڢe}��\qZL���9��Yخ&�#Gq&��i2ƍ�9Z�R�Q���hP�G �v�xq�� |%ӛ��H������8��	y,��B��z�|ʲ>�>:�h�E����u�ɲ��B}�T��s�8R�z�A5$�o�mc ����W�{�\҆�M6bW�O�mB��Ijt�(����w����X��5�ҧ�M �D�0�)!M\���p�`D�:�D��7���:y!}i~��.8�f�Y�y�L"�,w?
��r�M;"�8�|�p�Z�TX�T�j~E�F�.w��{���7H�Z'&����"k�d��E����!�	߄�R���`�6�H�C�ײބ��	�O�vNCXY��"�{XH��1j�JA�pU�1��%��D���#��;r<9>��l��<���8U��r?��QJ��BHc��� C�hJT�[
#�2�����^�z�[�[g��(�/�ljU�
��
�"�'3���i�)��Q�3�ͺ�]2jH��S��L'�A�C{�2��=���L "����Ȧ��d��pK�����i�Y����Q�&���6��o�b�*㲷+�Qs�=YԫU���O5Yo�ezf���7�_��_@m�X}��/��U��.	�������KK��L�?�Z�P̝>19\ƭo�閮��^> �_~K�D��M�N�U�=�}E���}��0��E!�$C��ג��Y�/��n�&R�:�g����L°�t +�0#Rh���.����'��㗮s��?��J�?$~�`�>fj�� �8�z��{œRRk�J�.~��ã�A��}<Z�G��wl���r�����|�B�k>�(�H�jW7k/s�M5��G�Թ(i,�⌑@���J�S�M�*�]�n� �c��m�m^��������\��F��h*p3f�q�=��s�~�٫�;	�8"1��@�?
$
��S<���b�6��T9g
3�����yy��\�hI�lׅ����z���<k%D�2m<4�J����F}Wc�
ؔ�.�����n�3Ź���g���a�,�蛠� g�U�a��8~P_}��V=��&�lN�,[�01�j�F~P�v��
�L��v3�֊��ݘ%9BR<�������l�"��s%̏,�^�S�?+���r��$��{�1�S����-�z�eC�CG:�yu�Yѻ�8�O
��F�sj������b��,.�fT�*�9�h8���<_r�s�a�d�v_��Lp�����SEc<:��{^)�(ڨ}z�P���e�>��u�sT�ᖀ��7��I[����H��>h�����F��:�Y!��mȖCC�K�`�,�O�d��c����\}�ׂ��,��#�-}{1$�����C���RY���e�}@p��=�R[`ZM�2ŵ��zf��nU�5@��J��ji�	�Î��+4)�$)�"O��Z�fD��T�E^Ͷ��+�i
9<(0T��ӷ�y��@���r��M]>/kQy���t_�t:��cYW-]B�O~J�j�r��K#l�������#|�e<u�?$���ژ�$ H0 m]J�ϵy���0��ɂ��q�_&��
��Dce\�*�'����o���lz8�q�)� �˨B!� ��C�2B��k��Q����O�CJ�9C6��|<u2Ey@i����k��$0/&��4z�P�L��E�����4E?��q�I�͠_B��|$�lm\*M���T���a3�ww��P�X�
�d�MaG0������D�����<A�ބ�tg"ѥe3q���As�5�h�n�|�	����Pm�޼�'�.[>� ��5������~G��y�	Ҫ��[ ^6r�Y%7��f�s�ÿ��=��[�:�q�E ݜ�9Mㅻɇ�o�#l 9x��~쬕o-lEʎ���;�&�������8�X6�w��0z:n2����I�'O�\��<��	���BWl!��Nt@R4\���m�Ɉ�D�������Bg�HI��qP�``��z��n�=�����B-sóS�Aa7��:8ND��h�k�^�3��>B�9<�pQwQ+}R�7J�m�|�3˼���)c̋���)&��Q5��N[7],� H�������Ӈ8cOs1y8�`1������>��V� 2��|#W�o���2F|2=+oR��_�^
7�F���;�$挣9��.L�X����}�=�P	L�c�y8���8\rt�bBUԷ�w�~�B�$x��UJ01��QD����Dm�$�CCl���XY�?��Q�����*�6TI��"d�ӸD$@2�m��1hZk��>l3�+p5#0m�Uu�tL���8@:�j~�U:B�&ݙ��TUO|\\|��K�,��k�m��p��m��ֈ�憣\q"�g�P�ͷ�y��;$�oR[ ��.Lc�uT]q3B���.�6��#z�6J�ܖl��� "�C��������9����d��D?m�:P"#�����3��1���4*���Du�2�wg ���}4k^���IC	�ő��y�e�_	�L�\9��c�H�� �X�T���қ�5H��h!ss�������r6"�0�d�HFK����@�O��7H��eG��i�&�F�j�E��U�!؇�D)b�{�p�;,�����O��S��4'���w�!z.��}һ�<m��	md/(�� �	����Ȼh3�7ėVj&���="����y=V���~����*q��ߛ�69&�������ҩ,+�s��=�wT� �?u\�S��f̍��U�{>M@Q>��y�dL7F�@+���&%g^|���AG�3��	�W�l� "M;<�=u�����T�.S,q�L���+R�l�:֋���(���*�ݠ]wXReod��YdYk�2b$¬>J��7#8�IG�,��I�Ґ_���^姁GRQY�K�d?�X�}�x�"��7�� !�	��d�`��'����ު�2P�,�u��a�$��_�����}w������2b��A�|I��v����%�Fj�>�2�X����Y�\�(g0�1�	a��T��d�ֽ�IH-�9*�Qu���'-p��B]fav������v�����Q��57f�*7I��;L����dc��b�#B�2��z�:�3KpL��@����}�e�Wg�ow�p4�:��-��;-��̩�AF����D]e���UO�J�iȟ�.#�bF�����|���|Mt)�:`������v������P���鏀s�s�]Q���·�eNd��X����q[��d�p��)�k� ͈�g���F��_y5����HU��0�#6���AC:��nH�#!����Њz#��J����K����pT@8��AX|���pX	��wМ�C�!pv�g�7\z�_�!9�`�)o�bWJM���~�LU^��RÜT���d�����E��YM��|~�ۚ=�WC�2y��߀��s�ߝ�̜e7��ʐ��I�xn(oa�6���f}f��=���*�t������[���&�O�M^��vK�����|7O.
f�f���80�j����Qv$o�ʃs��0�"��)�����䊜W��?y#1�ρٹ�h=zy�?L�*m��A߹Ӫ����c���7B��V
\E��ހ��2%�MJ�=��(|���p�����n|?�4��c���Lh٭9n����
���sk�/\��#�)�Г.7�nQ��8J��3+ 5��8 "��/�w���R����<=�(��WDjMOboѲ��{h��8h� ����G�ż5���Y�!fc(��MJ�����Фm�l�d�{~�>#	�e����{�&��7��Q].����'8�M%���[�w�ǀC�f�y���y�o��4�u"�Գ���0��C��:d\V�͛t��o�\��{o-���Z������0�4S2��f���-F�4�g9���������:��X�fL���t[q�3˺���m���������ё�,��8�P9�S��@!w���Z�H08<��]����܊8��<��!% n��FO;�C0�N�ȥ2Il����7J�=
�YdbQ����d

t�D4����I��Q�=j5�M:7��u����)e��Vܔh����7�#�sN���Y|�FS��*�xQ���nL����$�a�/&���LV��oGSy
�g���e�(F^��A���.#�h�x�ڡ�bF �����x��!PV]���3G En�o-�c��-5�H}�Z�9!��L���P��2��h�������{M8���CD0K��÷��.�R���b����R��G���s���������(n�1��T8\���Խ2Np��*�Q1'β�i�_��;߶b���T��U	g�jW)�o)�N)�6�F/y��h+bl������o���f�-���z��N���u�Q��vt��
I����F:2K��^���9�o]G�q/����%;�6&NG�g�'����"�s���'J/����G�)���KC
;��ޅ���3|ǡD���R>y>:,go��t�$� �Vw�Z�W25(9�Cc�'`e��ۻLãP�Y6ܺq<�U����Gbg���4�rF6���\�e^���Drۻ�,l�쎢ت���ω2����)'��Q9
�O��:"�^Ò�pBU�&���wgf2=��C��=��C���9���a���݅����m<[#��ǕT���WDͫY���_JH����,o�Z�8ޒ�_�Ŝ�7k(�����D7P�I٥�}	H˰>��Y��'��v�rR���:�{���m���ST�G�Bs��fc�W�.��Ť�k(�h��sK��+�ѭ���>V:���':MO2 ��O�Al_M�l�$1�u�$5o�����c8��S >;=�c벖���hT+3\o�5���L��K�11�W�(���~�X��9�Qej�.�E4W��4G~���,�z�w����z��RPc�*�L8���	l�}�?�W�VvX��kRh6���DB���ar��,��f>Q+���;P��#0'���'dP�M��(����0�gfy�ۆ���p��p��k�Yo ��PE���J��R5�4�"���.��Gh�!E��VU��<'[0�K����|-�X��?��W8�m).s�u�GT���������؃�T˜�Ʃ���Knщ�Gj�ͅa�}�~h®�]�� e];��4��Y��:�4ȸj���O@S��-7+��b2��z��ōj"\F�Fe3D�=z�KhR��V�F�PC��8|)c
A�*�Ã�pW6���]�V d�%�|���D�g�O�y�"��f8yr1��*p-��������H={���㔅�Oh �M����_o=o��HW�^Bf�vi���VXZF

S4fh�J�f�s��	�����v��Q7$	�"�L,�_}�rd~u��֤Zb����r�Qxf��ZTsLK���0�\��e��PWFd9�T�E����m��2���eЄ����b��3��$�i&�uAhS���Q�8B��X_
�Dz���B���tB�"�PF9tIh-$�nc����&w�B�#�N�v�e����9¾�c�t��^fv6=�c�
6�?Mܘ��;,��B-�_Iv�_��)T��
T�	��n�G��;��,=��3g�s+>�	�7�*%%���D2��0��'~��K�;ُ��)6r�3ߕ˩��'���R�-Ӂ�I��_��]�ciઃ bʇ�a�٦Q�C8��l�G53�a���aFIңTE��/��as!��5gU�f&��M	ϯ��Gb%k�v��#iG�C��W���M�u�J�%u3�{����)�=�4�Yx?E𿭘��Hl�3`g�7�{ܝ
��.�N.Oʚ7Ye��P!���SÖl�Zo�9�\Ѣ~�CNT�kǹBQ�ԩ)�]���J��W+CH��Q�f܂͹�ڏ����ﰓ�4|��$��`}�~�W��r�W-�6q�|��U��ab`5�,Ik�u���e_���Y�o�k�>W�yh������.�hi6Vy��jA�]/���T��@�[�
�7#R�1(�QC�3��`��l������5����߰�(�>����x�y:�ð�V��4�~��������1��R��[�e]�ؕ�z$#{S�OF��{D~G�'����$�)�S�������Kq(����fс�4�ܩ��: ���>��Ġ�14��t=h��N�3�yfCM�Oo|:�)�Y�j�Յ��� ۫t����G�����eM�<ߗt�/���$D���w�#�2'#�� ����q/�/����i1� ny�@b.�"�.��,��z�I���ÔN��$"?>t����p�ֽv_�a���`n5T�y]*}��3A��u.�2)ʣ�m��>�=?�X9����/��e-þ�eP��)t�y$�-�OLgQ�,T���!�۬=u�|�u��X�ڙ*�%;��M�A]�{�t36Į����9`�ўX��1�EZU��D�Q�?��!Ic�h��B�����\��w��`�Â�HY��<���M��q�I	HI�{M�1[�$�N鞭�V�*��T�
�(�o�[��'�G%��Ø�R��"9-�@��Q�l��T��5��G�_:`D��`��:t� ��o';���|��.�%-�՗�p�V'����8�(���0Q�sV��c����4N�ez�tQ�n \�%������eC7*M)9�E{)�ߓ�M���B%����I�2��a�_Y��'0hT��r�*��?�<��Љ�i�reĶS�I�3@�V�2��v�����u��c�+��U��i�[�KGp��E�� 񹁟1�˂�?��`y����K�ےp,�M��+�����W��65����)�Ƥ\������[ڬC��G����FA�礽�U�_[Mj4�R�UT~4���z:���v��`-?Y�hl�+fAt�"�닖X����%&H�%.�an֨G�a�ٴ�4�\Y>0&N��c�H��"/b�1.n֖+�>ܶk�ƿ"����/��{_l~����@-3��%O�[s�d�� ��A����MӄA�?�&�����]�z!��.NE�$���=��_�d �峪4�U��C�c�����S%X�p�����a��1�>�,�K�`�@�D��B�L����QG֟Ь<]&mys��2*�8vW�	�5Sْ�8�$:w�X�3�{��^b�32�L�y�`f�X�Jz��z�7���v���c0����d�h��X�{������}bn(��\KI`���m�x�چ��e
k�P���5�%�F��T�6Ub��R� �(�F�@3e���/�g.`��g-x��"�UI�r�-��{�7��.�ɢ���0R,���7�z�O �(|���"�����o��1t��c���/[��+��Z#N2���.����%\��sJ����;��Q�Zϝ@�w�®��C��<H����n�.�
�� ��D<�eo�nB��gtI߬�-�G%6�+.�s�Ҝ�D���	�喭���:��m.��0wL�xP#��:y�F~�0���\��-�� �^�Yn������!�)���* ��ޯ���b��6�O��Nj�ç%
<ӧ�7W�w"O�φ��L*!3[�I�}/����P�/��Y��5EWu��JX�A8\�a�.`�&���o�b��ț�rX�](E ����������'�*�2Ǧ�xd��$\�T���i�%�v�=4e_h�����Xk#B�h��\������7��c�Ӟ�:����S�)D�;j�f�� �CQV�CC1�<V̈́��^q���} ����pO�٬��#~�!p:*�*w�&����N�Wn����@muuI��� OEU���Z)�
��.���P��� Ϗ��;�8�MkH�|�r��w�"���z?�k -HHo-?^�;f�|�E��捝dHCX��$4duwKF;��<���Ø�q5��
���EkS?�@i! N�3;݄A"N$��y7�����o��p ���9w��	�1����s�<�ԧ%�fM*~����xW�&��+v̦���d�� E�&��:�U(�9��,���/���;-]!z��K�BFS�P���Ov���1��!�Z�p�C]o�E���Tw����]P�Ar�!�������-�x �f����F}:�Z�y��5�PmV��j�H�4�-�$HIf�6j�b�������z\o�?����q�����HMEƂ��Sb�m"���ct�dr���?��P���C�7�r�ⴳ�p|�~?��@�kH���mW݄�P% ��'��ʣT�`�]�W�������q=���q���O�>��.,/#�
Pw~[GA���X�B�mB�7�	�5Ύ"�$d�Hk?����?]�s��ϖ��79K�ejy+��(=#__U�=}��w�1�6D�,��Z����P��|ǒ�mf����E)xY��b��d�Ӹ���W��Z�0	C��\)���Y��O�N���]p�s��	�O�f�i�vZ��* 16�#��	���
�u�� b;(�V����p�g��B֑�p!�]�֨Y��"~:�����l:��ItIg�E|��1��2
�Ĉ����V��q}�&�@yJ�=�1�K�1�Ɔ��N'�3�z����H��8y��V�SS��P�"?'�	s�����ukI�*a��Rs77 �����W5%�K��g�hy)q��.#6�]ۺ55_�}ݦ�jE��n6Q�m��&��_��zTol 6zc״MM��l�)Ԁ�D�ݻ0b���Q#/V�ZXsL�罷i�V|��� gn�3B\�z<OYրD*�C���L�/VA���
��n5P�V�cs�X���O��s�6��N҉s��Kge��������92z������[$q(�]���#��ǵ���\h�ydQ����~�C����.l�����7��e�6"�F����Uo�I95ּ�_԰|<<<����$���~[B=No0�|�ǔF���X�O[4��q�:��{�F+$;R΂�n��~~IKI�Kn�k�:�sc`}U�5(��nY-����@�G򑢇�ʭ��̜Uȼ]���n�h�̎�1�s�=f�fs+���
;�����,�]u������r�j%�:X9A�G!}�s�x��A�ЛV��q�{녘ƾsC:'��_�M�?m�^�}����{��̫K�"J�y�2����!��N&�������n����z-Z`�
��^8?T�X6K�[nla�����3�,��Ux+ޟ��1�_�H�D� ��l��K��d��P�o�;���gAP��]�6/�j�Z�2iu�����w��1:��+ד�I{T��R��5��0�U�t�T�k'\f#�Ì|�l�Ԗ��z����4�-��o��#�	Gᆞ�x��� sֺ��G-d���x[ڠZ'�&>Ӈ�����+
���kb>�'����Y�%��Yn�hH���ް9%�ۍg�c�Ä��$O�+�,Y��hO��Üz]���dy^(f���s�6�`S+@��#m���K�0�e�Q�,�.�w�5 tu/�w�/T��Y����w�Ԥv��p��{"*����OV;۩���$�?i���!����x��$��n:Ű�O��-�����ʅ���r�A��B��кp�U�U��1Dr2�Mҥ�,*( rް������:o�H·-:̺<^���Ё *R��v��ԩ�{�pac����"��&t��}�Op�M�:�:��]{�_o^�e�����P�_<�Z[/t��>$���%~�����^1%̠�d��0��C����2)��h��C�]ܜ'K ��,�=ȄK*;�.I�4jr�K��"�:���	�ʙ�����'w�����b=�����~��/��[�~����4k����H��Y��l�X͟��R�����{��Ƶ�"8�K�5a�s�c�KD�ծ����;l`1؉��$��e]��94]���FM����8>1Z��fk�sN9��@E�>�'-�e�X��̖7�v}<�I����ޓWm<ӳ�� ��%�����zd�A��j��J�^��(=��_6�y��<����x��5^����t=*��֪k\]D�B�l�e����q����Ҋ
B�91�MW�YO���)�)���+�&�O�7�B��u�|MuHNr5^�C�xk��c��W�:���"�6�gu͊�ܸ+e�V����n���Y��ለ���j�S�R�j����~�fI�ܫڃw���-�A����`��'���f�P��nV{K�{?�f�@��*���& 5�;�((�r�� ���v�ʞr���(�6��p�B�Y�qQn�-��=�@���u�ɾZn�?h�ϵU�_yڬ 3 l����קhn�<:f�g�O��P(��& �ƋSϔ��tz�9%��ԅ���#A��YV��V����[�#qn�
���l#�,����a�B�E���$��5�uz�ϰ��
�[����C���ʊ�/��q��ө�2�'*��/���FxX1��Z{:�ӡ�3�f���ĳ!�(D��]jx��9��୿�pN�g�]����F�Kv��vՍ*(\���EB�_�~�ϸ*��yG�q�9�S�m�����!�0o�<,q�_��B���:��d�>%u|)���(��l4���!E!�}ZB%����k(��AL����n�8tV0�e�me��px16�Z����k�;��d��f�c�f��$LMZ�mŏo����F !�;��++F;G���o\��8~���$Ȉ8�Um�+��(�^j@����,[���AkV�l��nN�K.��PF X� �0����y*�-J5����S�+��:�)fҮ>}�"�����A>d���*�D�{�Y;K!����9���$6����k.)"?~�'�2�3�B&��VO�n�!��K�N|$���Uţ�r7F�_�L�QΒW,�٣� �a�TԽH�s�Qr���3�ܛ�/������	�X=~T�����Uk�ޅ��^Ԅ�6��}.7U����j�Ys�G�'n�y�� �2��`\j9���ᚗ.�L�Gc�)�z�{G
�`~p1��٢&	�Q!���x�id>�\&ǡ/>��NDil��+e��Y-�	P-&UЕ��[d;�f�sL
Q��~ ��c�0Ā�%��L��������ڣ��l+���PuV�G (Q�.�k�d\�	FZj��ĚN�1J5o;A�!��Wg�F���[�<mS(�;Mq�Dw'oo'�$��6�ք?śWv������[��E�B7��]�3��bu������r!��<�����j=�>ދ��m����xC�.�_��?7���NZy���X�yU�Zj�K�I��p�9��4>�T��N�ϲ��!�z�3�i�;9T/�E?S�Ѻ-R���f�w��Ш�K���\�P���8���������Y��2��V���y�$O|Ԃ��ñ�V_plN�f�1�c������,Ch��c+(4u�����&9�B-��G`n��I ��m//�Z
2��{��}�Q`�	�X�ei����0�u�c��I���8��tn f�tvX	 l�o�m.�?�z�^�H4�hZ��RJಮ��Kٶ�L��V�s��<9��B�����#�s�a#r� ��{�ހii*�H (�O>���fz��R��5X�ά��>����:��%{�no�]s�Czp�w�(n���nۅ�c����L;o���H5UO��#D�i6n�8|67rYa�~f� ���a��F�0�g�b�5��M�	+ݭc�?���,�-c�~3c0�%�-T�����.6�-?����bp'��'��F��oQ4�_#e�񏏾�5K���$�x��}Y]�C=HN�	;��FY�����p4��u�uUȕ�_\�Y��KZ]��FWt2�f��ZBt�=��|�J^�(`�s�4f
6����/ջ� ���]輳N-t�f����}>w+�z9)��������yu�@�~%���V�������F�wt��*�o����}����(���j���hzfG;���(8f��9����sߞA*WJe�ɟrG��5�P�=t_h�_V96�gd"B�ӈ��
��]핰V�1�-�� Jh��ʞe��$�6���ĥ�4��ѸdYl�;��~�!����Z�*�"���V�.b5�D�EeW.%��%�7���ᲠYs��O��ʫ5�I��R)�zL�%��w�7��|������D�=�|5�k��}O�茶-e�C�B1Sq�\������=����'�΢_��9�����b�YW�41^T���ծ�����:ˎ;�:���o3��f=�e�ܷc��[�\k� ư�f̑�X]�Y�G>0�~DB�"b� 9��]%��]�$�uir�p�p/��ŐN�G:��Wҳ�Ĝt��҅��ߧ��������.9p�Tx�:�(;%աq�u�C����q��
hwrp�j޼*q��1�a~t���{�J�ߥ����nD�65���9
��#���9�g��)f{ܧ�w��J�9S���d-*�ba�l<�v��-�\�e� Mў]��@E�>��D��!�{e�U2HN��5,E���D\yH	��g��P;U�}Ts� ��uR��("T
��g�)',�Zh�����4��8�27���6e�}��[��?5d�F,'_c��/�#�QO�? �̱|)���7� �D�����p7n�3qrMB"`��BT��3�����
���*�����/��;ˋ��M�]��K)v��tz�~���\�H��B���Z3&\��og�X�˺��3AP�Vb���#�Q�l�ť��70�<�ړ��i�	����Ɔ��
�F��g;���YS)�����%�3��=l�P^ph�xw��YLn)(k� tM�����>?���"b_{wO��h��+kF�>Jxu�8To��'�Rwb( M�ϲ��S�M�+���7Z�Ϫ�*�'�$)&�o/
{�Kk�Q��P^�v����%i$ �= EO�����=���fE��^/�Dӯ��?��tԣ�zMᝁ`#�C<�S
_A�-�1���-MX�a6�
o�����&υ9EJӛ�����6��$�eS���(�[�Y�VB���ƭ��wC?�k��]��IR1)�vc6=#��T�j]�F�a�_o�Kۆ��ٹ�)�Y4�i��d��y�e�c�@���5m�Hqw��%�T�4x��2N�G��{j��o�:5e�+�-q*ms�y' X)!!qj/�8Cx\���{
��WIv(�m�>��~��T�7��<�D�]��!��b��i@��$�v/tN���k�.��K�7v���/nQ"��B'��7�Lĳ���=��(��lRT��iiJ`e_p���3�E=�D1����3���5���R��+�'z<�'�ۘn^�"a��4&��i��N4ݚ�Y��gb�E�ջy�@]d�G?n<�κ��Ow�;��I�`�f��ts]��b���;;b�p���cU������!3��>���U����7wkh3Tr���Lkv2ǁ��r�b\ ��b�@�(�7��3
��V�ONa"'p2s��i6#�C�s(pn�
���t��i��kz=�Ä��	v�����y��%�<~�F�𓁥��<� �1� a��+�C���	(������i��{m�+	�c*����CaԊ��c� P��� �[=��;Pj�Z%?þf��5Ih6D�'�~؄Zbܛ1{7��md@O����&�q��׎3y�ӟ��I�I��k�=��}[�2�5���C9��.��m�*yW�ÝNw�a��9%��]���@�(�޳�p��7�SS-`i�_B�u��F�}�f�#^Bz(�,�s�_ߑ�#�<�#�6�Ŀ|M��~5	πVu��A0Z!2�GYjUXkB.U�|!e�m�i�)x��9Ӑ��`�0��!�S�Mq�A {6�������L>��o�b�����kӂ�CU�Bܽ񱊉L�m`U��uw�\�u�_i}���
S��s]� 0P�C�=K�@��w
��!׉qb�o@���!Օ��@���@s��)]V� ��u��Ї!|A��SA��{s{�^z���<�;>��b'/︶�Q*�j7n=z���8�dt�L�FW�R���@&3��v�o����<d;�Ѷ��	������K�t��1d͞��d�D̮��{����̽�
P��z�w^����x�~'�ɜ�xN0
�QAU[����
.�C���ÿ���F��(����w��[�]z�%�J/h��ȍ6���Iq���76Z_H��nՙ��c�δ�$%A��20�b���?�!�I��b"%T���
�cSy��D5��dղ�r��X��m��-�cB=m��+�P�_�>ynKhk�N���l�mMx`%c�����3������c�:�5�F�"j~��`>��!hqӊ�E@�<җ�ԎQ��%"WM٫\���p,��D�ݎ��e��95&L����kכ�A�#aYa����S �����ۅ|R�Ѯm��d�Z��؝ob
A�����̦_����f_��{���.!��?��D����ZȆp�w��h�Pop���#�_��v�x$}��/�Os��T�C�r�&�}=��&*�N���#���� [}&;�8�v������-Yf/��w��M�jm�2Mj<�L��ߤp��+�}w�
��y��U�Ύ�2�:M�;LUX��ʩ�PE�D)5@�����kS�?lqrD�!�Ȣ*v[I���o0�t�6 ␹FG�*��o�ё��S��$���N\K'S���G�55�?zУ�A������� �z��Kc��I�%R�*s5�I�˸Jl�^�� �?J�Ɣ�P��`R����]�� ���"k�o*�m��R�Pu��L72��
3�Am/���m�PM���Ĉa{����q��DHc�sRMB��T�ϞB�Ӿ�Sw4wst[ ����/��@A����:�"b�Ű����|�i��s�$����\�.�e�+t�F��;3*�ќ�j���4-�{&:%XHռiP��t��B ���i �M@r�S:{5�������ɤ�@�P&�$>��H	�ĺS��F�}陏9u�:<�����#yi:Q-�@[Vb�ㇱ�����0�s���K�L�M�K;)������3�vϨ���Dq��lyؕꌎV�'�ɅL0<7��I�GG����c����3C붕�E����/��?����jKE�*ooI*B�I�.����A�Y��N?Z�_s^�<�2�P6C�;��w:�gӍ� �dl�=n�P�:=���3�$��곣��U�-���Ex��-�,/�'{x��¦���l�Bi�4б�t�ɣf��p��ӄ�\� ���ފ��⾌�oKxNo��kZ;P�����l+O͒�����_�ɭP��$1��gZ�@܉����2���mКR�ip�� �].uI��.k���Z~lr������w�s[��퉸#>i���
��=S��S$?E���(&Cx��U&~M
+��Np��j��>3�Mo�'@�t���,��]u��g\#_Q_b����BƤ��<3�P�`��ӧ����0�:�ynӛ�����pQ�����C���<zӘ�6�C�æ�Rf��A�E�hO�	{��P���*,9���po����~���U�	�*h��*B-�$�]�D[©T����%d�%v�+D����m��(@YC�J��la��.��\~�b#�a;��|�Vڅ�n�K�6�*���O��_��_}��x�F�e�$+UvE��SM��0W�����m�-��F �렃��A_o]��Up��y�t7�,�=���~�7(u����jl7(s<�Rq��`�/n�����o8�ڝ�������)����gp�7q`B�+�����ď���oxg�#�v/���?��ag� 
��@|�[��˦P��.oCsZ�_��T2�%ϡz:>1���L3[8������l��e�:4��>��a?u��;��Ei�W�dZ��
ު������+kb2����'�%����v��T��J)F���=�'�m'㬅x�ķ��O��3o��eg���QG���y*�6OoK9�ߺ��QڂMg���8��H��2���ӿ�Y��8�;\�3�p�5Ɯ8����k�qඓ:��M�`�b&��ɉ+.�EAo��["x�<ˍ�K��*e)���0�����
�0��dp F����*�W/y���l���F���%��V#�Ӷ
>����Jj���-�\�_��vq���Q���c4�o ����fbӂډ^��PʦsX)�uN�7MVE��`�TƝ����WTa���YXQ�0-���v�� x�s"hA���������=h�'���
��p>ΕR<��UBx����D�!Vge�5j�d�ƣ@�b������+��pI�eq�I��lo�h�߿)��]���iq���Ok �XB�'�&(��dmK\���P�/��(-B��������uC�.5� @'mmc��yH �׫�8J�|�,���/'���$�4;CD�/ �yY#�.�B�����y����IGb��\���
��BV�
Xj�樥���9b�%< ��Dj�/����]����27H�w��e�s�"��;m�o�@K&��:<7ࣲy���𓰅@�05�e/C�b�ʡ~G�||�*D��Ֆ�����CrS���r�eL C�͐&a-����.�
��L�˭<�m>��c�}q�Y�%8�g��0�;�����E����zy�qY�F���FƓO0��g��t�Ug�n�ۛ8�K�A��Q<?Usv��7�EVI��d6o��I���"��.�,��W��a�=��_��j�\t�(7��M����3%��;Y ��k���0�B
,utˏ{�	�~ ���~9S��:���ȟ]��!@��OJJ-{��G��=ޥL *�ص?D3G8�d�]J��N����[	]��\qUUa�ۅ�)DY�g�=TG��%����)��jL����������tP���O�B���!9e ғ�/�ۓ=IO%e-����X�3�����`했+M���O�-�QPi��3�I5����þJT�
��O0��@��.�/ʌZ�g8����^��wS �ȷvЁ�@�1 {�w04��S�g�O�4��q�Qp���l�3�j$v�İ�T�_F�DC�J�xXl$���9�-�I:����s+�)/���*r:'���H��t(�7��{@�T��رs+qzU��q©��`��\���W�Yc)3��L.���0$~��N��*��b�=�H��!v]N��
j�|Ջ�ӗ�b��h氄o}m��*����@����jl����� 2's�]��&�l(}��تTU������a>7�4c�:f���KQ�k�ܜ)�h˭�����	\Vi������H��
cc�uEd�+?���]4b�������=줿�Ym������vm��*��f��T��A��[�w�'BYe����B�SYRSg[�iMX�s��J>�|٨τ�xo�V1�K��؉��[��K�H\wc���I�ً���<6(&,��5��Z�b�eD����HYl	�ayx�H��z�{P�����J���ݒ�����B�Dw�8Ũ9L��>���#>HFg�Y���e��^r>Px'����u� 	&H���/r�B��DV��g��8��[,�6v���[I)I�2I߶��Wq�N{�����2�Mg��4�a�v�r��=Mf��7|��M`:�N�G��lE9��p�$H����)V�Pn'B�$���)'8���,�r :?��gBʋo`�L�QY�5A���g���ֻ��f��>��Z�X�l�[�_m~���Ǿq&( [����}���k<�����:�x=���Br�L�-1��y�|��D�x���m����#+�լ6�gvA�[��!a� A}���J(tL:$\�
Dμ;�2�;P�M�J`$�����/�w�	.@�4�v�D�%��x���4:l$q?�����w�/�M�J]7�}J`�`_�F�p��-1�/���_�_���rb���ɢ�j��x	q�2l��'ZQ'��K1	�ěՠL�憇F
��d�<C�.�u$g�%�g��C@'��7ts@C^P�0��ב�T��ԇ/yx�O�[K�(7Im_�D�An���3�Ê�?nD�`�[�~7h��������u\�L����9�joעԤÜҏ1�5�t�9��6�Ȓ�2ӎaI�%�Obg�z�(�C��=�ƻ3n;
�:�0�Ly����� ��`wk�҈Zia5nj�vh
�B��[��Z�_z�����g�nԡPl�P��p�m�7y�`#�&��#w��{<{tW��Ȯ ^"����h�8E7Rè��n���o��o�u��VB�dp�lv	��Jf��M��֖2h1B��C�1�eҊ�o��ј�$��,#���K8���6��t�o u����s�Tw]��C�F��^��ݣ�0�\<ch3�k��̱Z��F�5���WI����`��\�/':/�l@����>��L�%Y�m~��s�\`��VI��873*�φ���RX��+����K#2���"�,3\AqX}[�r�@+�����|�&K����$�;\��w(Y�*V}�b�&�Xv]�jД�y�(diz�3�����[ꩁ� ��v.�ش��w��S���
a��M�U�Iٱ��A��e�]�L���G�������w�+U�_D���Y���e��Њ�g�C���n<��7"`|����\��Mv�'��h;Vo�SWb�����MO�eW��Ya~��C~�������d|0'i���\�m��>�&���(���}��Q��G#��Q��%�W
>	���/:�q��ס�[�c��>�I��u����3(F��`���S�lT-����l�q�H�\X�U�P��F�0���PM��c�)��p�A�!���tx�'Z�R������g=���R(�5^׋q����f:���N�׃���fZ��5�U���MX�wP���"ڽ�U�\����������%�;�������������>G@�1��Y��=K�o!/�[C�ř��<��BY����Z�
[����z/���V*���OE��w<߄�+D���ot�`Eq����4nq}}LPе]*'����b.[�0�tٰy��-�D3���xĳ@~�+$�lȕZ��q���O t��U�*����A`��������Y���%�RGb!�@f�(~��N��C64^���?�$1���+yHw{�o:��r����$ �T�^���˒n����ѿB����w�^8�����$�����ĝj3=wy��k��m$snk_�I���G���\y��?h����
��=�J3�~��X���Tl�� BÐ,��M:6>�4{{ҋ���51`��V+�)ZE�.����:�_ll����5�@Ű��>���	�u��í�\6�'[�8	�4�I��$$�<�ˍ��@����R>�#eN��Az�^�`����qy\��^(i4�$z��������$;�����'J�C\_#^��I�o���B׎�WP�c��W��L�kZ:d)�[!��B.���]O���4������x-���q���hl_K�A�*ƌT��Z������~���1(գ�|�u���6�"2�U���h[�Z9  ḩ���{���oȡ%7���aqQ�{�1�N����3s��i�H��#m�&�v�/���´Y����TS��%�
�y���6=p:�
�j&���y#�T�-P����6���	:d�$[���;�!��vG������H��KZ����/�t��j����]���'MLS�`���M��]��&§p�?�1�Mq������b\���]u�ۡ�	�E�הGZZ��P���6MY*^�m�&��7K�M� ��b 2����0��mE�&���C��i\�bT������0���O��I����z��H�ԙ�P�:��"@sá"��sPi��I��&P$=��֪��'��:�:'�r��$1����4�e����T�kH'�
푫n���x�"O@�Dz�	S|�#�?tT�8�V�c�p�%{��tm�� �:��@�%I������j�@`�~�rJJb�11�`Ti�b���$Qm�|�=��#��Ӻ:�-$OT!��?���J���r���e�̉T
K��5����кV�g�T:8�gK嶄0���я7�|���5w�q�u��%4��<�!�[���6�{�3��w[�VQ����e�:�V� R7w��? 
����	�+}\|7~G�� ,U5x��`$���2`�sV�XaH��$`T���I���v��o�`�)��g�Hx��YA)��x�Պ,��_B8�`^,�~�?<���/���� ͛]�*�[�H͌E���Z�kkU�d{�C�q3��[Ghr�;<�5J,�<�a�Y=��^z���h� ���� �P��]}�O֪�x��0��LBi�'�x��7�J]P"���L�]���V�KkRs�Cgu1o@�{�B�wPP�kj<��5#=;��t�b� ���1�>��2�Rtp�N�305�a5�m�����1[�:=A��^%Y%�ݳ_vWo��+�<3�ac��O����m��\n�>0�i�~ݪ�c:!� �b!����9��s�w��	����w�1Z=�^vT��� �Y!~*0,]@w�؟�ؽ��B��vޭ� NtBq�)�J�x�#r�g��~W��8� z��'�?�m��^;��'�ow���|���5��nI��La'r�Y��5�!���֙Z�6^�>�/�bL<dо+�p�`[;2� �a��^0�Y S�/�v��i��J�� �=h���4ڵ�NT���`���q@X�Ȉu\�J,�v�������~���kP�Me���xO��;]!+61Ճt:��*]=���&�`)|۷�lڛf���"���	z!�@,s��_�<�ML�:�kZ1hR?"#CȨ!���V��O2F�+T�5���.��C�߁م��㧚���Rzia��#�7В�������Y�8��zHn�'��;>��k�����ߓ�p���ċ�jl�>ϲ4Ϳp�H�nQu����|<����)�W��Wzt�T�lOڮ���oW�]���#T���`���^u"�c	����0��a�N���	R7��Mq�t���9<蹘��n��[���X�'�8�*ߏjٶ�pV�Mxg�u��4�:h7�Jg7��N{z�ι�(��ѰThS<�pW�Tb�� �"3ሮas	�m����J��{-U+���Z�����f(����t	��+��AZUZt|0��Cps�.@ˋi-4�V%D��Ȫ�ǐ���o��^,�����t/t�ąg-q�?gǺ%MO,��1삋���N��\����������z�;��o�N�����;_�D� �WV�+Th [ŏ���@�x��ןƧ�� ��;��c�p�zNd��^hH3��a p�m��.-f�D�{����B�>U�.΍�W�ڡߔȦq����)VI��싶�˧���U��9&�Z��1���V�Ŭasޙ~�ֽ112���M�������q �=�;�Ld��U��[���J�t��	����?�mT�'�q�f���}�y�����5�SR��L�t�*d�F�9S�7,�CM���|NA��$F���W{�3,�g ����?���a	���d�(]ւ�,g���`j����7r�6�/���:��/��	R�0��d���cV�ڇ����q�X��2&��#/��t��5�a��\"3�}g���L���	���a�p�KA��Vut;�;!B�w�t)v<��<X�F�]��j[mr��==���3W(�.�ނ����8�Sm�[X��<lP��<���W�Y�&�r��z��"������ׯ_l4��e��A�/��Pe�Ն!,]���?:�N�w���P�Ԛ�d.Z�d��`���UD���	xHM�c���߉��UG�i��b8��
C�m]������Q��2|��\�M��,��l?
�T:��I�?�g�^�^���w`��r/��h��!)�j��М�D���� )�n\#�k����<OD �:��X��oO*���:)(��h�j��~CN�ӎ��`�;Ut�����r"�~�j��P:�������:pA�6��4�����u��9���2qA���� 4��W�G��)NPM#p��զwDo��(���a�%��۽j�!O��� $��Xޔ�|�J}�E��8q�"l��Ō`��:s,��R(PYr����q�N�orhR���`��ɘ�jm�)��:ް�����|Jd���Mfp�ӫ<#�v$�7��"�p����8�s+��Xo��ig*��q�A,��N+p�V���P/f�iؿ��rc�%�q��=��2��W5fe?�整�Y�_5�9wt����Մ|ix��1d�꩎��(�,D8yMG �B�g�o�#�\r���:�=�[�ʚ2��VU���2��1������x)�_�(��!s��Ht�h	�В�h�^i�-B"�](�f���� a:��lk��~g`j9%�����O���&w6����
��<X����P�#�	(�r~���Qd��*5`�;��w;�c�`s���ϗ���U1��b��P���ʻ�.�N���Vu�T������uX����E�B�S_&�0~�A��rK��|���p��	��@�#����B�3����`D>��5�%7�l�<V�q�Ȏ����p7�mOq	$'}w���U�u��_���?���S�>T?���	L��t���dn�����Q)؟�g�]�=�8��#7���k���*�t�¥ҿLJPv5.�Rk[��Դ�3��;���i|��kYb���'lsIm�@ P��л�)���� c�<5��W��9�1�X}���x����x˛NA8��R;�Ɖ���UD[F�T��
�U8}%�Տ�,��y��w7ˮ�_�H�����v&e)Ì�n����
)��9nf�S���ҝ	�X�!��8��SS���Bf����6ҡ�{Q��r}��p�Z�0="�^�ϸ��V�MEษ���S�C�J��E�R�l$����L
:ɕ+�<+[��<GTڹ!����<�3D����n�ce�=|~��9>�j�>c���E���
LVMޫrQ��^� y~$�s�|
��B�F�� �#_���ة�?�G�.\�Y���0�9� v�]g���!
1�;�*(�g��X�v�b�9�� -��Ɛ�@Ey�!�O�Fm�9��,_+w��cTL�[�+�ז���u�Q��
�C��dq+�^z����<���۵��v��U�Q�aY�v����D)��qF5)=$��$q���܊�5�2�(�K�bo��� ��Բ�I�~�/ʾ�Q�c(��v�D(S�Z��V7�椶�<�a�Gŏ���П�=�׊L}+�f D=��e�a���;�~d�ݴ#!�Xn��`	RK�TLP�
�/����9#X|5dy�4��l0��t����4�%a <�S���~�_���Ô;�,�!l��xh�� �Ś�Tl���և�L��Ͷ4�l�3�.t�7����Ǽp�r��8��d�qCS����ˆ�QV�O������o�0ػ��[�|;��"��gR����J����+L�⷗]�./>óg�^���D��,�*��
w�5�+��9и��\��7��N�	B/�-0|�+��F��0�L��9�-O:E��
~��g�踵�� y#��"AU�����;ȿu��ٌ�޸�¯�Z�>\Hq���0����'�:��<'�5`�2���W�wѰ�<r�k�����:!IL���N� 1����v�m�gŧh6ue���P`g�2����+v+��ªK�R�� ��@���X�Y�#���ԚR����3���fa��Tmb~]�V�YB�J4y
g?�tj�Rk3�2[P�S���Q4��0"�64��d���S�Fb�Nw���fICљµ�N��*���S�m����2u��j�o�1���.�ܣ�0��:@��N���k��|��缠M��ͻ@����r���Te�4i;r	~:�������xKa�i�̋N<�U+�ɀV�������ը:�ZV�<סGȗe��`�\(�u��y�[$��}�pi9�l�}��Qxp�t�r����K��d'������`�.�W8��S_�P�CU����2��8��}Ͽ�J۲��>U+����X7i�AB�E�W���v��4�RVn�����]E�w(^��v�,��\�\w�/~��c��*0Q��%\���p��Y+��s�����H�^"�,��B~jjєw��<��y��W}���0ۋ���EebP­�Y�)ˍ�A�ggh����Eٌ�u��"r�|��Y���٭ًH�67�g�pFw��n���z��m��������i�g�(��e+R.(�R���4�2�,�;koΩ@Κ��S�Ftm��_{;���}Bz�,@�%��ѵ�{+v�
��O�A��r�o���r�i.:ϗ��W�tu��2����2ft�`x{�ӌm{�4v)}:b��aD�C��R����^�0@�?��)���B���W����C+KvC0j�zS6-����V�i�Z2��+�$n�*�9�U�6��(ײʖ;/�/0���a����% "�`M!�����rP���(=��bܹ�����2���ˀ��on�Zc��v���&>ab��J��%�F>�T����n
Ѭ�[���h^@C�B�����vg���TR��� Lq��W*��D6ofVD X�6��j��r�[(�j����׳{K��E<���?N{�y:L6I��^n(<�?�.�-�F+� �^��{B#��4g�!4��/����0����s��EӡΡ\[��x�~�vN&�V=��H9;�AxBc���ԅb1�nJh~�8�멟_��.��<>4T5/���\1��r�t�"l��l�#o׾�5E�}A=�3$��dy�'p�:2Xi�-R_�&�n� �������[�I70���������e� ��C�qձi�,dr�>�9{�2� ���=[JR_�1��E���DlaX������,�>��M5|��Ma�޼�|O4*l�����[v}8H�����?C���@�ʜ�F���?M�bY���+̾	g�qQ��.�xҫmenCh&\��8q-�6��Y�u���� Y8���	Qh�i���˂h�)2��d��������,-,
��߽�я�M8���w���>x������%����������+X�t�C12@>��#@<ݺ�v�o9�͹�LG�W����gI����f3kV�p!󁊴�zo�F���.[�K��I�6:%��e�q�w9��2X�@0b*�*a�a��=`�!��!J�"gn��lr�y)�P�8�C���7��w�����������0H��8�'P���[�-�x�1�.�F�	!{)R,�g�$a�z]�;$3�Io�� K��ϩ��JX��Q������g�|�y��l{ޜf��tq�L�R{hl�_s߸���EP����t�/�4��a���6�$�{4t��҄p�˝֢�<���kcEr��"}*LӴ\ه�6ܴ�ȿ�syC4�oSy�r����vC2�I�^ щ#?��ׄ-�/;�=���AHQU��h�]M;�q��C1H����:���5h���}���Mu��]jM������l�~߃TY��t��/'^�Eq3����Ѣ��"U�ߎ����b�t���&��a𺆖. u�r8�s����DT��GHx(�ӄ<��x�&�����ڥ�_p��4�=�2��z)�o���"�Ņ�����$��VX[��BlQ`�"Vِ�'��k��S.�F���g�]�pܼ��F���	.�����,4��%����V5�yVz�I�e����s㼪����,*9�:�דA9y	��}�UjO!E�H�M�%d��D�u���pn\y|�� �\�R��R/J+fK�N��7���ä��{_Rl��_=R����i��P��Q��=�u�f����T{��;	WoyFCq�X�'HK9��k��WO�M�:��E)q=�:��0;��]�đS��G���ˀ(f��v��I������tk�eO~�=��z����u�5���8�4���$ic��F�l*�	Jj�\Ū-�Ӎ�2�u3�d�� ����2�z�ؠ[dM4����4`��xd�=>���Ʒ��4)r9��!�k����{��J�JY��!!���0�Ѯ�Ej�j_>�����/�Tm�O}��&I�w����1�0_:���V�|6�v=`��=籌����ﶞ�����ps}�⍽f��G'R6�X�=+�*����h��I��#נ��owQ���5r	�I��)��HrK��_��k��6�P���$;��mAe�-�̓��?��1����iq��-@ ���a\���v ��[|�_�Hu"�1r���R��3���f2���}@�Ԋ��r�Ms�ɢ�iZ���w~G�+C+
S"��2���g�Uzx��\���Mلx��Z��Cړ�����}?εЌ�1K�
�����}/��?
�]Fs�O��%SH �:���bJ��A.�P��oF�8�' �'�RG�G������'E��w�Lf�vWv�В!%��28m�F�3�����G�t}]cY�U�'��*����Yi�u�_)��_���g����t�7��AG��BI[��_ET��-Y���}Ԭ0��<	��RLJjo��k����)��̊�)o�YH����b��L7������1;��Y�3$Н|5�P�Ru'oe����<���ʷ_�k��F���&+,u�	tWܩ�ʃ�j���
��Cg�Tn�Ղ�k�cK�У�}�We�鎥��!�	w�|���Y��$J��^8\F�x[�*<A�u�Ȑ�N�|��ݱ�`(����~�P���F�����$�6��`(��ZՒ�֦�0��RIa��u��:���j&��{�S'����c`(��M'����nҐ0؟�'���Ԙ_o�ʹ1)��^(��q"�H ��Ko�]q[-f�F�T���8���T�F�8�-Pm�,"�A����C���1���mеe\�������#��,�$�Y>}K��؋�b�嘮8_��ѝ)��U�S�g�����7��
{�a�ᷛ����熰�����y�|�?3�Y?^��\	�H���3e��Hj����?�<�T{�y6�����|Z�	V2`>��`���'��`3�4�K}ٍ^���I�^��,6��9��[��������[�輣���̫�$������>� {�m�+�HgH*�{����J��N�⇆5�|��G��<odT�5gp�3a�s�����ap�8�K*����/�=�l$[�
(��;)崯+^
x�a1KRE��M��}�%��<31��y�*Ñ��y�sne�T��χ�|[���k�w����$�VL�^~���kHF �X�wIa5�L�TP���;��~t��mĘP����w�)EQ�M��	�!.������Xtг&��Q��� �^��]�z���*hD�2�YS�~������$S��i��G��~��׳[�7��tB�nn"��]���%���@�X�E�b�K)d�~�����h�$=�%�.0Oٰ�u? 暺����,k�K^�I����O�� �� ʂ��%ۤ�v>�nr3osx߷�n��}W�y<ɇ�âu�R���,�Riq�H�`��Wh��ڨ-��B�{;o���&��`��D�D�e��1���ZsY�s�v����Ydw���V�T��C���6w��!K���GG���^_�>ҒR�M������a����V������v��0v��5W�U���y5sk��z|�
�!�*A�������@�����,zX���b��0M�
I>�&L��Y���P�j/�eOzC ����g+Wd\��wO�q�u����Ϩ���J���M�H���i��&��w�s��;M5v�m�Ư��ZC�n�j�CPE��IB�h�TK�}��L���)$ß �ͫf�{ J��T%�C�2;?a�vA�f�Yc=t���\��]�j<��0�Q����|!u�p{l��� ��'�E��H �]�3�&�. ���i��♉_�rsWr��ڿw<��>�HK�$��Iv��6�Ñ샄�J``S��D��}�4�ƼR�[�M��?t���v�C�y���8Vb��jP��m��?t��IИ�w5��ܿ8�~Ut*�D_M����g�`��L����*��A�A��Q�o�Y�]��j���t����C˾���J7�7��� ��m�M�b��BW���Z��)|�.�����TU�В�{���o_K��10Jw�g�641�$W��?�`�g�����28'� �k��A�
��W��Q����G�����r�������̨j���8?!N��HC��a��1�ɬ���L�7�`���ܟ`q)6q�<���M���z젃��?����/3�X�ɾNF��9e<�K��yDZ?�n�;s�G64eB0�?n5O�7�	��܅5��6��-L�_.G1#�ݜps8ss�1��?cW��AW`@��N#��e�
ZYH4������P��T���ȓ�@��A
Z���&���	�ay���	8BM���
�r��AnC�O�0w������q;�R��+D~��.�L͏��ƚ��P^M�4���KLI�%�"��ѽ|�F3� p�8!B�z�N�1o��;�qnZ��՞"��]t�6DY�t�������:�	����UI7���񊋯z":N��es8��72G�Rp���y����*k�U�����(-��D�.���49�ٱ�:|�& V��q��_.
Q�g���&��5)	���4|]ɹm]�]�`����C��ZX"��hn������.)ܐGiS�N��9��""�K@�*~dx"��'̽���7��NS)ER|��3�1#'�Xk'�W����JQ��Ύ2����>��z`�A,��J�����9�h�����1� ��k�����*���5R��o�:���y����C���ܗ���,�!(?��X�pk����0�Kvd�oe��n�=��G����ĭd�x4��˿PM���t+DѦ�mi�k��*[��~KJ���t#����y6p�vl��7+�D��� [P���Q �4� Y~L��T��(Ȑ�)��4����^��~�&�Dh����a=�6�گ�ky�{��z=i�֙T�v�>�e14��	��!�5��3�Sy�_w��f�$���h�Dʴ��7%< �*�Pz*�t^�c��mڴ�Aʷ�x�\�RW+{m-S�c�{�E,�G0*$M�v��T����z�2&lx�5���^���%G2c?@^)�|ċ�q h�|�5��Ȟ�<�h�%/uҬJ$U��o q_�/��r&oqu��k!�R{��8X�ym�6�ґ���`(l[�:��T;J?�ǵ���@[q�E��Zg/��o���4�?���������d�(4`��� �l0�;d�̆^�(�� �qX���$p�~����<ˡ>j��xд.�:�:@��4�ػ�P�T��E)�7�B�AJ/%�ެ�����3?��x��˿�?�����&�~_A��f���]z.(�qG�Ӻ�>�;QC�#Gj��$���;B��;�3���0��,cܠ���2q"V\�Ժ(ELPK�l�F��|1v��NC�����$HJDI���OXNe�I�uXL������=>sl%�0y�г�H���^��T	MpnH�c��|4�\xcp��~��d��vDK`��.N���WP^�c<q��_<�����"J���~��T�nGb�Bvfk��'�;��G���$.��3T���j��^��'4ѫ�3�����B��U��p+%ʘ�fm�kkL
��C��:e  ��r(�wҊў�q�W�]@��I��h�D��Aٕ�K׆Ă���V"�u��As�E��	g��nn\��]鹑�F������ٯP�8f�G��a~W
>e��]J�;�4���Պ|k�>JC�� ��>YI���bx���Q4a�+� D"̇16N�?�^�e[�6U|4�Q�a�OϋA�$�!rr}.Q�<�o%��x!�E'�?���"�3.�&ت���A5}�n/O�����Y�����5��f��LXذl�'w��WNt7=��eF�ϵ ��� &�}B��Pvs"��W����u�d)����0�d^T���"�%��'�%�g�>�k:�S��.⾡E���y:?H�}�Ќ`�;U���@��G+dU;?
���8s5���!!r:�-��D�����'P��y�'O�u}=eIW����� �#͖�V�~a�����K��3[��� ���+�e�I)fꂧ��)��IO~
�/���Q۴"��xb*�|ԭ�Y8��}T��$h��0)�Y rA��n�,�	���HX��$kM���:��ߵ�H69�r�j�c=�Ӷ��.ll���Z�Q�}��#�Y'3I��ы��;���Z���D���("6S,ҫ�k�M&�giP2`	��p�4o��:��c�cx��Ƣa���N�\��t�Z�k�F�D>��:� r���'ޏ1+�ê�|LU���%)�����y��A�k�p��r��Uj}P4A)�ȅ���:��QCK��=y�b>�\3����7��"��v/-���Q�qp�/��-��PM9��ܬ��"�Ma�|��$�_���T}��tpl�27����4YQs�ww� ����S�-��^o�O6�2s�xLJK�/3��p�S����鮭*��������#P��g��e�7^����}��7��
U�8��Ynl���"{ЅW�Q����y�q�~��� )��.��Z��8ne� �X����ф��B���v����)�4��`�d���c��]��)�kEU5��+q�R�s��t��f5f� o"<c9�Sd#]�|���{�*^n������Wc\4W,w�q�}�K�D�
o�X#?�]� ��K��=����z/G�p�Z4~�����|��d׶ŵퟧ�Ӯ� ��NE7	TI��}*�1�˶I�N>	���Pe�����No��f���Z�0�V�:��5O+`���|��B�k��j���TkSɰV�a#9��5]�s8
��O6�@�b�˫c�C�{3�Je�~�����$�n��k��ZF�Dhf1�L�c�)a=S
V�k�� ]��<י��%c��?c����V��NK�cz"j<�k҅��ܼ+�/�:8���L[�@�&'�G���*G�m�!�9fT�מ����AR�N�`'�ǁ���)S������ Y9%�1D��~T#��3���a�VVn	G�G��<�b�����_	���1���y5X��\ZU���yoG2$�XE���7���Bu���ҠP�[{&&��Wĵ��YO���	W�C'QG6qyϜ�C�����<xC߰#��b(�?�ͱ�\� ESꄟyo�[I34u��f�cW%�Tg�G�V0~�}N�r��k��[�AG��/z=k�(�4�s:+�%aE%��d�����
v��@�YqR���Q�%���[Xcs>�~މ��=���Q���~>��wT�Fas��a�陘c��e$JpL�R��c�}+��P6��$E�U�R1�����2�%��qs�fp(7�ʞOahᥳP���|-��ǟ*��]��
��ee������W�7]�u��i;x+ܠ��n�#������K�&�2?�DI(h�t��\��V�i�l��-���h�g�z�w�����`?9�Uٙ	�)|���G��TT>:��UjKK*��	�8�Z�e����e�/��I�p_V*L�zZ��Q�<b7��ļ�Rٰ��JY;�?qe8W��4�Ϡ���Mi��b0#�r���`�ʩ��%1M\�l"S)�-^�"��_�iHqɭ6��?I���@�$a|0S5��b���Z�O=���O�*���f�F���!h?"|�9;���7f�r��ڮ���ղ�U�tQv�cmN�
��*�6<.8���p�$�~�z����ayP�/�9��g7q�<���5r�@��j�p	�)t�*���б���9��l����hx�躮Κ��fCb��A�m�s�)}�crY�������)�'�#b�k_�8wވ������ȹo^��p;8��`�'��l��{6qȗy��H�|�0���H�#��G�i�<���W��WE'� ��)ԯZ�|}��*C֕�6�����l��f�"�w&�����l����a��[��Y�J7R�wE§�+����~M+�cF�0�4̬������ʲx�ŗ	�T}�{H�Bc�_�,���]ڏ�%�#�r����4=$s>j_�^��8�w@��݊�i��V�r۩�~u.��5Y���#���+�P����w�
�p*?G�h���*���u�]�Dj�	�Y~M�U5*�1GG(ٱMJ�?���մt/+��aOF��T���+�/�����W�@�$b� ��!$R��I|�A��,5۴s�%2m�:��8����F����XgR&�b������[(D����&�p�iV������܋��H�q�ψg
&�j�M	X�n.��t��ぶ���ҥtFo�Ч\��*ҭ���Y�,��"lQo�Mԝ�,��KU��U�s�������3,���8�e�3��r�Nv������U=�=�Ɯ*��OnMP;fb54(�-X=!LTq���Oj��p3�#�8q� �Z�G��b�oZ�������oa�݇$x2���*��<����m�0��_�8��,�����1L��R�Ǐ��4��0��������H�
j�c�{3*�X^,d�;i���W`v��Lq
�_��n����6K-��x���(�c�<!Ń�ySD�*���ےf�m���p,�}&�G��B��WI �������F��Y▁|z�;�p��W5j�W����H��u'�Kb�����X�X*��*P� B�3���*%	�l���y�O�������%PgЉ�֚Rޜ���G̼C����
�q�Hlƌ�k���Ӂ���c���(9�s�c�^ӦքU%$�ÔO��I���|�"(４�|�>벯:~�q��Y�[R�>��.�Q��,�*
W_�YYQge++|7�B��ф4F��69�Ae�8���,���V�ڥ�p��4��˝��	]��fr&8���#����ݿaԋP^�qu��*�2�3J�#y��C{��c̿��~D8��a�<7���[�jr1��J����٫�r>����{VЈ#��QI|����s�7Aӱ(!=����ޡ���<� �f��}��*�ӽ�4Y�m�6�|wNu����x��pZ)���V�`t��6(������L$\��z�	/|f���l�݋M�u%D�i����̔��gp�ׇ���F�&�#��G#�?7��l�T�e����7m^p�/m�R�d�L��c�_�<�v���Q\���'��}�鯀Y��bq[W��q�/*Wd�\�q�EɪMֆ�+.J���O�LmxԵ G��0�'V�
xyZ�ؖ���~����u�Y���Zm�Ǔ�O�!a�mz�B<� $ ����T'N�E$Z�,�t�QqZS�J��T��~`��p��\ٺ�>��Y�0��f�0�U��>�p!��S ]����y��9�Ԯ����ňp�S��*g�Aa�k��mYtg�A��ˈ&�N�%�A��RA��a;/=�3�D!�>�?���[��Hۊ��-LK����P�߼*�)͐���Y�;/8Ѵ'���.�r؈�f��><zffGD힢)RsS��-s_��_����Rz�U۷�-A~��|cKQ����~��O��`P��f�33fI'������y��q����6�@�ǲp��a���7[)n�pZ	�&����]?��չ�Yk�`ی�_�՗� h*���Ihi������䦈W�t%&��c�6Fʈ�a�(�JF4 ���2��d1i!|2�)d�R�
Kr�6�=`�����(e���f毛��he@!q���ݾX�������ܸ����6<r���Z�RU���zB�^��3i�~��B�m<o��z��Su��"
�KPY��ȭ?��8�BCՂ�JKIJ�x��46`�M��/�����^�@b�^��E�p�3֭�0��L�כ8�>��m��_�a{Ή��$���Y�R��!��49�v��8��/�ߥ�|����]��8ĔΡO^�H6t�F�)�4❑֡Y!>����rp'2�����ud�bf���>q�}�=���X�tI�Jܕ�"��٢����ڂh	&�'H�Ġ������;'L�۞�Ϲ���	�k-f��*9dH�P<�t�wtoE�.I&�K$�oX{ϘU�J�_��f�(��������0����o�Py�Yx����֔z}�Yn�4��M���/[���b������<3�\���ONFp�A�׽��.Km�f���l ��6�2�� �jXk @gy	hx�@�N@G����Ы��V^S����%5�/W�Rm�x�V�d� �omљi�����ɼ�,�:ɰ��"�O��筠dmes���#�C1x�Kc�,u)�
s�5h)t���+�UU1�#4	q�a��dĶ}���;e��oޖ�8?�58��o����0�-h�����s�Ҁv(�GW᪞"1\ON�EF��W[[���� �% b��P_ y�B Dm����z~�#0�1U_�wQN�a�����Y�xs+�^A��Y>9/j�%�f��v�?�YT�C�5.�>�-�����	�+�@=3o��v"<+x��ݟ<�L� R�-
�p�1�H��e��=������!K]+��\��}rz8�):;�^�8��i�<�0�E�@�s���*nV0et�֚ ��\���qt5�.�Ta%������z�sZ]$�[�𛿬��lBhr��1��Ag���>����-aqT�W�0�/a�gB�î��zi\���{�'�ک�+?���i	oM#%�Ы�P�B�gĤЖ���wR֡���Nܪx�nK���T�?o���f����r���W�s
,��Nb;\/Ð��%{�vu�A KGy%%��@F �'W(6[1t(y���E���fԾ?�l��0���xe�m8>�
������ׇ����:Y8�
W�b*�U2}eLwm�0�@���st�h�XsN;����Gˉ���	��̏qk�]=��v�˪ˬ�~�W��	����$�8��4nC���w��&p]V=����?F ��� �Z��O�s�v������1$\K�i�����O���ǩ�0�kA�]J�����5/���ԟ>���6y���8�e3R���B|�������&�@����j#Q���TKڣ� ǯ�$��W4�� ���n?�������e��!�q;��Q����#�J��^��O�rB�y�����6"Q�.��b۵o0����� ���P���p=�����Qةw-���}��#@�1tu�Ɓ�3�8u0��*�