��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7���_R����7aPN���BƉG(SѴYۏ~�Y3+�<�&�L������ḍ*���u�6ᓜ?j��{|b-ْ�(��
�����m��<�B>_�$Y�73�^w3ՂR{RC�OS%�$I� m�X�n��0ucj��K��r�˫�}STa�����yy_�]F�3�ڹ�m�nt֦ ���aZmgD���g���J�� C�vr���^�7q��=����xݭʷH"-�"�?���x�OȺV�6\2�0(�3�!o޾���>A��z�k*�p�cG�-Y1q����Ѧ��1.i���7��I-'��?
�_��lg�g�mV}�C����x�c��z�ڜ}Qf�7�i�7�8�߽´'�5~� ���J�Tޞ��oj� ��>�	Qn�M=��s�@k�`W�(��}��l?�J��o�6�}��y�V���n�<�RH��>bk♶`p�ڼ�N��T�WԭH�=ؙ%s�w��,�a&�]�����ms)��kѲ7	�U|&������P��9/�l#F��Խc����5[��Ƭ��5Ju?� 5��Ǎc�E/��u=k�Ï��`�����4�x�d@��69E���>�~��=�H^�p��qII$ ��_B_��D�<+^��
�0���H��S�\r~���D�%Q8ش�[_b�E�$��zr�52�ù��
�LhY�4�ઙ	�=�E���S���6F�?v,"�Fח�]'-0"5ŎYab��R����c
��/Y,�_l�S8�R4W����Un�P��ƁK�7��xo��8��Ce���妔�X'�k���t�'P2�F���_���!�;��k��ɋU>����4���� �v����q�b=GKgc�fϮ�_�3ʾ�5\�4�&;x�]���E? ��Z'��J��$�b�h�ò�m|����ë�y�� �rI?��O�\��%˥t�@��62|@H����G�U�G�g�ʿC�E�q���R-?{��0����Bm��^_�R�������w�׫��z�~s�YA�ۂ�-Q�u�h2R~��h�qȂ��߾��m1�������PUp�i��Ir��B���X2����G~�\d��M2�S�yǅ����zˠt�;��cV(��@Ԫ�q�����c.mI�L3���g�'+�� \;҃myd˕kO�>����6�Q4ibt����չ�Ԓ��i�62�!7���^��L|���~͂�k	� 
�=[��{��t�����a���E�8u�=��74���M�K�*�e���R�a16�hM�B�դ�n�Fx�ɿ���z#sb뱰@M5���%����w��+�5�ف:��I����N��:�oO1\�Z�.����(�2E�w�ua���'D`5�D�}@H8�֥m$ʻAzȓ>�I4�g��L0 ]�TA��-���9��s�p  �0C0��U��%����2r~!{�*� K���K��[�aU,���UR��id�F�2��sQ�JJd���� ��x=
3���LQ�}U��6��GC�ug���8��3Nm\�l��g�⇬�Jf>�ڄy`_�A]|xt�D�U��!���Fyj�F8�ɯ��25�Z��o���0CZ���P��pX�ke�m�o��N�`	 RR?�Ram�b7Mvs���(��UK(�*A_�:.~�O�u���&�6j�t�%�wMT�ʤ'o1���vI�t�^����$�;E�*!+�b#�+8� #6�'�Nt��W�����t�K��p1���	�aˈ�~�?я��ګ��:�Fg�-O`5@T�߼q�F�P�Ra�}K�v�-���K䶀�-���!�0iB��ʅ�h�����Qޔ���ũ�-C�)�_�A JFU��c�����Ws�1��{����_��R-FТ��o��	Rd�B�=ި��;�Ҷ�z�H�1��!�2�i}�ow%��<bh�sǣ�,�(��!<�y���9���J�`��A����c<7	>����L{�|�j�/�8p�"�tng�c�־���b��1�C�`8�~���-?9mX�k�wT�b!����y���Y	� �t~��3�������^�j>_"�����r�dхPMb	�e��������U��;X�S�@)g���~l/���ѥ^|����3ʨ*_��}�|��N0�q(��fW�W�r�#NC�C�I����A(IS"
X���db�����