-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
llx0gQ3/NvTZIc1XfYPgNMLVsMGbjUpMs6W4iXMYhyEtCMfmsVf3eSGCjAvyx2UwHoDlBnUZIi8w
JHOOIZb4KYGOpI4sZPR9N/4ew0S6GaILR9HilRKi59evqwuOiMdw3F74Z/R6sJscWyY+anfF1eNI
mvNaItrvQOmPfie77gv5yj+oiLTzJVrwvsduD+/Q2O4vGX8Gogb0+0cmbwFGr/NyMXTqDfD39oT+
Cyh5tKskmKrKXWs0y7FskSXIJLlGI2M7Nac9vUD9tsYMv1yaEiUnfecwRb2LmBMB2S7nkhwAVdns
eZq2RI+b1B8yOWnIY8xkXW9P8K7J04OkjndalQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 11888)
`protect data_block
3McaXyQw8YIJcZgp4Xeud7iVIYEKqh9h6ZOBzfUAaHGz83gQt5tOjTTp3uE38HK8jKqJlySYY8GJ
DpJQ86e36xvUpQVyninc6SraAaOiLkC0unUsnuCTVg8r4iT5RwqDbrbaTm+OehD32JgHE/17X/Pp
YhPIBW3f+usXQqHLF5NZ7IrWBQbG6JGZ5z8/gGI7siVoy2geM4b2JCtfBhndhDyIJktjvObjGR9o
pQdsq988UxAHt1lCegVc30f3WPzlRqm3AY53Uo32eKgWOLk6nMOhP0VhAaA3g2K1LScD/F8Hk7Bn
OIV79p+kwo17RHPno6TTal45e+XdCN+tiob5EwLyQ8GapA2Rti62XbTf4IAXS5EFnodgY/mWey9I
zrmll5NQu+kSpdMNPBJmryOf8Z9LkHif9EqiiwUU08RH6pFdBOHEpLkKF8XrS6iAkHWBHAK6+Gn2
g0dP4xOcum1y7qDjDMZwQZ/tpLiCuZ16ZUVHvW2bUg5dfKXNNVkIp3IuUnd00b/asuo60lGcYhVT
4CgBeKkwKHTPpGBiQ+2RY3vuFEwxdrrnmDDDuMH4tk9xJ6RUBYbYSeFkx3vJH9YwdAYiAKaDPT4l
kzpcgqYf0Btu6FgxG3qRS87zu51Je6mWUM9/WbWi2FNBTPT0rrV1RoIiF8D5eHdSIT6/E/Zi/y2V
+EvqPAXkyPLMincRkZnZmPKSVQ5bq9AzONej+/kPLKRYjwmHHm9K57yCwfinwO5wN9SjJqIOndHC
ZHWTNaN6iuWS3gxWTgXU2Z8lQrRmVjzqraZiOUE0HgHpwU3pOcfozNOewXtz8JCGRIu37z/hch0X
Mmg2sOUfEjKF4mknzWkwDLQAp9yEViH4+5m6BDV8d3kmQCl68BiLkCWRaZMWTEtgB3cJtb6/K8J5
wl7F5FlUCgFfdc6J8JQuH+75HgledH3xDxRsarkW8LMyuD7UejWg7t1f3yqJprEY6rZlZDM6EHTK
5DC9pnvyYsfSJIewTuoljqNV7JrkktZU9qKKZXJ4clSt/UCTcRIPiA1acE5uZtk4HH9Utt1KkTEV
YJzzUI4YTtr7rzdEZM5MQiEAwxYHlY0ni4CrdyVJ+BCPn67Q3tiiTEftpRg7mUgdz4Y9nAvvHzrT
i3wXkSo/novnh8htLkPo1a/RRtq3M2I+SCEVFdcU+gX1Yj0pXQlVwiD6ypCRtIaKON+O2zkAIyTI
px8VYDrR49jA2Yw4Oiy7scWKA+XDwVrX6igfp5AQZz1TU6io8bOHxN4DGmjJwcE6yj9pjdDubdEm
BBqlWmHqrE3QEITfKj0xzUcIz93DqfQxZffJ3v6ovixyy3NDtF9NhTAttTKa98I5FXwju6nBFQYq
NokdRwlkajtyC7ZNtVvlmlhuQk39y1/EMb/RyZI3r7aco6VmYuFuQsJTeBkprl+B1YEIcRkYEOIJ
QHKBzMthRRjEquBVD+w4z8xt5afAmh0b2m2vTglEGAS3VIHmEtKIdeR/zWKwJ7ei55P4lc9ZpOMa
Kg4F+M1Js59f8Qmezdk6fXMupLOmJwuo3y97JmqKEI00NZc27zGc2RHRByXXXaR+ndda5Dtgz5ld
4ex7sb82xWKqP/kxmK4B5LML4yk2a4Ivmi4luwgqHmtRTO/Zk5GiS97i+uJzGYoVVFCsY8JswSpF
JbxMbULVo9ZaNIu/PsIGPneGJFFCYeC8eb+B8K8zwTNZ95u4EI0KqPF3oY/cmn4E8xQuzRtqMyKK
aP7TyC7dVrTrl6LEMcjOGF1AAzvbBz2ZXEElMK30u57Ai6/ro5Gv/ewG+RPMF9RlHBxDF1vdgkhQ
LEZDb4s5FBt0x9BV0n5TVOEuiiQlqYct02H0XEvMKeRvjFmAkT/ZnzB0Ek53usaNlky8WpOxQT3d
Z+xrnQkteBOfxJP7+gjubN9lXy3/rxaRoZzEtErZPU1Gr+aJ0Qdr5odP7gGKwUdfst48OiySJCaR
lB+aU9T1/82HdfBKpf4Y+mOPnQ23Hh34o282+y2RfOphyYl4oaOVmv6Hq0dP9KT/R3bK+S4WBnYl
3vhAuZ6JYtPrlBLNShjcsaP+uNq3Aq+K1oUAkj/uwmcPhZPtawsWbG0B9B570kKJDNs3AStbxSHR
T8MYg22s9sY1CIeiYrwSN/f5OoXsX2bwoj/PyaP/cOcsQinZ8bXx8RJEgmDooljWXODxYRCP6I4j
IuJELnmBXbxeOpMT0CBtLuwvqHZpyYVGYvP6/2VtoMcrvLZJlti200t+43Zx2VdRLsuH7ScHMo6y
c+DaQOGQbPiveIauE3YojQo10eQd8J293zCQwoV38OxcSPsfRorBzUGCd8VJfFrIMT9uBU71xAru
Fhb8xZoEH/HMCQcaMtO94gn4NKWhkrS0Gh2FcA97bBnzVAYdsPttjNmPX9PSgy4rSkTxF5TURyRj
oJ0h7bN0nXnCSND5QXA2po0sWg4SMG29DLqPulwUB4ls5Tg7xxf6RDzxRogZ3VFO0PvPYN4kgdVL
Q5jIhCQI9QgRrYDW9kFfAg+lqc6IF4tDBxTNSQQniQgzuek4NnXncUVF1W6OqEVCa53GTv+YKyVJ
0EqFDVgC2PXfcYwtBlLSKPGfcvtllcsoJXblJ8zPqewXy01WtvgmF3X/xPJC5mzdE5gqZBflYgb6
IJJLK8FDuF/S7eelVrVa62aOrp3MkVlPl0dyX5741ZlUH9WU+QsLqDslVYPXDDEsU5LbHs6Ncvp5
vuYCLpR2UieFtyl8DHZ+NLbNjWmukz1Oy3n0H5m/W/iBSIv4kNly/7zG7WkTK2tUG09obg3InVjg
BsAJrEFYeMRBSB/ZtBrGieubtvXS+wPyRTi+6/rvDikrA9NpybTXTzmcjoo6VGjDDY9GZQYkbps7
smbEavGOtSOXjcPcEQWqhkvF2VF6qzKZNSLCpIe8lC9XaSFQGFdRcWLc/x18RaK/KOXZ39aWRFAr
VQS9fvBqNbZH5RMYfJ5fBNlmodrRGblc+lolpk6x7b5bkkRKRHwjHvY1X0SoaDuDLQqfnWMiFo1z
3Z+62PFlg2MtM7yPwbUdD+qHHKD4oOmyavpho0n3HLhG6Ytn/0PM/QXa719ygBZdLAAx76Oc/it0
SxejtLqoZTOTvz99QHT000r9dA6JyL540x8SZp6SGHYmY0HxfRDEVDwDeH4Bme96GLUXZJT9LKPj
olkWibMwh4JFjew5MNsz3SxdwBRfZ4b23CFgieniepoc4UlM8Q92lE8DLtxeQxqJpii02MZkcWPa
YAZlTOXuBm8AszLzgV95YgNZULufG4y6pC3+ltH1NSrkc74n5DiaTNhCA9T9Hi/1r0e3xMtYVH2X
+I/RzWbiyfpufX7mu+dV1Uv3b/Gs2PmF8Dj/gYZ6eDG6yDQF63NIoq66f31GqAOvpTeWbmmo71+B
uYIbG36JBVROYkaEBnbQza7ZlsKcTKpJaa2YWZ1mQB9ExyQhH7Pn/43Rtxv54epM/m0RJBee4eyA
qboYorUXoCwNV317larZyTtsLDCw7Gzk8TrwFHpE+n13g8O3n3y3A+OVg4uqwRKXAKxiRSZ5CVXK
XNnYm3RnLoC3kMHudEo+79fgIFS4QkMvoS31HINwJXBit/c8Z4mdFyCs6HRHI6+nrIj4KKHBbP80
H0cQz0n7lTEZxvpM3IA4ZFdY2OrEoQmYR51EbH8tyLicbjpWevQfFNUtA+sk/vdpjAWZ0nmc0l+3
wCFbOfnDlQuirEH4Hbb/MCsT1F/tOESR5RnkDMTDxqf/sE1tkh2SI2afF9u+k22OqUl6EC1z067C
azlBOan6c7qJf60dCyQfdOlozGudfbMwIvC8Zxg5G9SqMWmfkNuovsXgaTQPDnQIJM+/0Mq+6nLW
Mtqp9NBMeTm9lz9L0iDoXBkNwHasjfswXuJUgHxvW4fzvG0KBEgzehwkJvSZSnHTiM0myJ12e793
j4cYfAGNzlVdABG2lRWU7MuDNlitiRQCqVVY0qgAzj2Ve0nGgVhfkeMm+FzLOU4m2KfMdLb+WbiU
P/u31gXGMejnmVi9ufN4IxcRl+1dmHsGM/MaMw/YCjLMpCWdbpsnULDyC0QrayF7cUWm9vFNp3JZ
al34QUrvJhb12v4IYihwuXti0lHOeKE5/WPyZUcn/PPzAwCHM7i77Fduoq5p+2s5DaeDX6ach8Z8
KDdcoGeWMLUvLakWh/5Lvck4GHAyr57AYBAM2B82rjPGVoeSZQgDSVXSrU2NusOe6WJQrKtkWek2
GQAlwTHY3DP+9I6x3oCutsC7VC3rUJ79YJlbRfapxvR4iWmugbZGxSgsiyLDK7WDBvmQRRIm+yGP
cthxRWfqT9f0QTi2Y8Rcj1vSHXRztwbPE7x40cEA2bwVX9ZKp4Ak1lrxH+ntj3RUJzG8brTJmOXN
swel8Z5GZu82QNIeXSai/WEXhSmRkGjtAKtG5fUSlx0rWJBcQJSF9OO/ykLpI0jR01B6zmcB19tZ
YzJGLX4lAAM/x8rRZWZXWr7n+sviy25lO/eqqj/kgX250cNAErHNFaczpT9yrKAT5ZGgTOChsTB2
de3sFZ4ePulUOnjTVfJkbT59s9wS3yieuFgHZ/CEogaQCQRQwxJvaNOQ7gg49iobNRtajVtT9iwM
gebs/DOrOdMjjVeek4oGsJ3CKcAkNe30qn+FzkeG9kqkzGYmI9xhoBRqkTghfp5rxwmIkXWuF4Ns
OyqKF3JaLLYAEtoKwo1a7U4iTjLr+pc+XcvOTaKwrejV6eEUNXtvjB0UTOJZqsxfPBVUfqb6GrEd
c+PaXq7MCX+JOPVnX0ju5Uh3TtFr/EGZkq+s5kA4naJtj5/ShchVWMwwbf43vPrsvZnaYqeiyHlt
QgkOkMvNeI3MvXKbC19LgEXGNEKIy++3VetOsH/E6z7AU6Ay0kMJKcavVrVqLeVqXT89v31fn6gI
K2yLOBEpI1akKeHsOr90gM5R4TOXJ7ynm8EyPNH5YzIkPY5ecrIv+rEDkLKNUU08uQOAyDOOgbZd
set+rNMKDGEXHbcS4EaiQhFECsoaju9Vz0aY7oUMttlRmhRQ8nhidIGw81fZ9G5ZN+x4U4cJpRew
y5Zt8cLIdkOXxDKS89uXXz947visP5SI6qpwVnq4dvVpK3CVFBncfzlaVTEyAH41xHhhmsFvHZJO
Rcs2ytVVmIEHIrxL0DoxWSYuc6lyII/2FqW2bqhw9LtHiz9GWbCnhHGExmLKz/KqvnYeYXBjDaPa
yP/uJ/p/rmNIAdTYB44iswQOA9TB4klDc7LwY7TA3PZzOxbfRpc6o/Qbuo6GireTqlxl8AREO4xE
JqbyIZyVGZi1WQMh6r67d6SkxJZfWNW4GM/KjcE8wc/8a+iKmsjVquioeu1LW7/1V3KVHLELHbM4
iVGgr1/QOZ1nugOkRJJgX1Z1/v4ZXQmrqNOQOkPSBuzPTGceHupKGh4YotPApDjby5R5hRIF4jNS
5cAc9Kg53n45N0P4axjBaOH4YHyabpASnEPpmnsVIA98bKufm7y+dFzaQsXR0UFonleySKjzjcku
y+wFmls5xretUOqp1B1lzXLHBbx93BqhKbTTsaBB1jsiuJSI4jiU/vyokEmYD/zRWTB4/7FGEJyi
qtc21j+bfxj+4m9DbUnZ69ftsFyRZULwXSJpeywoxE6i3jPZDegRyxNmLtsjrmqSHdks1goI+tmb
dKEYxRFZquo5Rl0flzlkdKRNUhIRRomlLmirHpnZhbdYcGk6b85vHi+35c7MsmJMQYnCTCjOD0oT
8Bb13EmDxcIPFfGM/6BZX6zFoW51FxU1lAL2IDtdNnAk3wscrnVSPlv2ffMZ0x0bSVjLuPmaxKry
IzxEOpdFcOrmnmtKs+jd+9bNnkziRwAHgbK3ICE8e51A109JnjLfw93VzNwsf3c5f7MLyC5h2FAR
ebDl5dHEmVfRrNn69W9OLmjUnn1wapMyvLjTJ0jkoQZxwmL9dywmm7bEFYVDRWDr2YlUgpNKfzyo
MBSO5YoTnpmDSV7/lQBlzGP1aYoz2+4SibEsi66EUxe2K0CbswnmSppT86I+bwHfdqxFsPFiLOvF
5sEjSnAkjjq8cXp/qNYABQ9GfKzaZFrpnn2I57fHSlqxq0LK73Jvct35s24nCFKVIBl/U01NXNPG
6prdmzpSmAZ36THRqejIN/26E5UDRoQ5Vj7PLQnhO8ZKlaXYpq7QtvBUDFxmc7RJJA6siAK6LvMe
JJSUwGSLOMeF2NjwbBmyub0n1QSqDQ7MaDj+aFSfOLofD7mC/+EFElNQRp1TC4pdNIXg24T2HiJl
38LY5w1yBSHQL4THOcqzTk5CwM0jRA8kocoYjFUu2Iyn2sExtVbl2R+r14uNyGAIlQkCm8YKMUes
8RlMuwTlAPm+KqzK+L69DRkNp7x7DuXcQ5Zjjn803hCZRbk2UUZkTwpIrELITmhRpLNoDUlXzYp8
RVdHRImYFugMhkf4Un3gEWofgSGMm6UMi92wOCRP0/olPYy+TXtK1j1kAtZL4BMK0XIxWboT08Hg
4E/hwUfm9ZFXq6eR7InO7THuQWerMClq5bZLPuKupSwKf+K/CxZBS4Z5Gn/8RfPbPR5CYq6DPkxp
WfxVqTXxjaepCDw0Afh5gzYLFeMcl+6U6QqQat4u+5LEb+4gSI1qhX28ngMgdOi5zJ28+ELfOmt/
s3l/xRSfrJFGHu5rwhy+yJv9ese7+QEJbAu+dJ67m4HSMjjse2x6U7ZS0UmOiwacKTgespsNTWHk
+hXX2xIcvT9Dmtgb7v1K2ssTrMuJW0tCzGNZZiSFO6+NR66iY3ldz2Og7UuoyE7e9tsfCesiFXHw
9X7XnDhbE3BpXEVfgj4fXsjw4fVfIMz19q2SvDe3VPahst3LURSWPqrruJtn/7cxLdTwrnYa4+Pb
fjWJxIDIs9H10gyBgFWcCJHFmYarAVjZal3z12o4l06G2mvy+z54MXjuqxEPWh9Bh8gQuwXUhJtY
ynkamGcLbCa0DUqFXj/1M8nO0mmD+OJhFrhkZw6KIMi0Uw1BBof+Tq6rKgLkngx8jPEp2FBA670O
9Bqw5DKWMQsWeX6Z5NVZ8LXUyheFKl7oZvG7Bh75zXq5ZKgGDPd1jCucRnQ/5gTj6zbYdThw3JU4
l52nNBEf2DKfoaD1Myt29ib5WwsylXV3KexYHtYG0jPejaFa6yAit07nd71rFfgW/DSjL3JzC1kM
UMcg9NmPZz3Oq/bFLDQr/n5BoVD3+hDhIwktamXqhPt4WeVOazSXqvPy/arpX0idrgmw3Qo0I9CV
kUDJkxsmXyurGazU5Hs9EWu2t0VlzjdH+4U3NyS5KWCGu02uoyAkNPwOZY7KZs7WbAIo7jxr+ZS6
mboi/bL5/5HQwhzqvfVoFixdT2wq6ilDBAXtXoDhGOR/z+8jsT2Bi17AZDsEYf/T7Q5no35n/do5
5iTwst9P+CqZfGwuqyf/hKYCi2Z/YY5cCL545NzfZ3VkicEYv4sP10SjaNS1gJns9aD5kzSq0ESf
1kDnsDIUtVQYgh4CqV090tQyrpE3gnRgsIxud5V8CHl6DfTuoIgTbshCg3hAmsDwfM6+yX/xUsob
zhlWHwwgXv1bNFeTvpyU2DKaCMlZD8Z9XpKca/QPvjW9v4vUHaIxu7MNJDXb1wm2pF4e7YoljjZp
QcAp7HXaxfYGCTE4QHkECVtTdJ8uJm9xWzgpTusD0ExUCTga5rQGvnuqkSThW6Wo8Uq1BjS24glN
+Hi2OX0X6QmwsuJ2ZRbUEpzP8LQTia8ffP/HnO1q5aiEbngdS21Hhs+t6zm5KZuLqUWF/SP9Nj23
ZDmu7pw7CCy+Y/WrwxWQuHt1z5uNFqGq7IS3TrbCDwp+ANYatHu9XQENywXe85k8rWVOSUseIlpP
c12JUsEpnoUylY+xw+Gg9Q7H9sARcaT1BwyrFp489yVGDrdC3iPJ2rpK9GI8T32cu1WCGI8CjDsl
iXyRn0x+L1BOPTr6hvH2So4qPsyctz+lgMUx86bw28OOsW+4gv3k0qcMWpgroZaE+eturAjnxpGJ
eEvsDjJp8IfUgvNvupgtdEOc7jrRGhagxhMQeGLONJEr8MmzofAtkXz3MufUcvL/h+pu3IqMU2b2
xboHlpQxWlbIA4CqBLygLfiuq15sfo0oCWbkf3JkjuNmINP7ou0YsVVqVye/2qRU04E/06xGpzFD
+7HOjiWlSx7j+SSXgqlKIDQHj3OpQCwPRyxISjATI8/lBNY7rA4IpMEfND08cnKcd9JHybeR6Fg5
iGpuGfhy4c2yV+0wbZVttNlwtQaOpqPfd8KTcW/TYCxTyL7ulahjM1VvzTN3QAHfvFcCnYIDLacA
SygSBQ9NM1Re+fgcdnEKIz+yz2rhhD6lhXU+1/xeZZWjNyCaIu3Mhvua7VVYBpo47fqmqOLVlVhA
jilYzoz+o8at3jnQtl0hQn0Yj0L7qq07gqcx5AvDMY7QvpkVEiud+IE+mR96yphsFpZOvMH8DE0v
EOfuy+N3BQ+AJlnV8Uys+E3uw3haatXyOKkG5H6VLVGoPYQV6aoA0ENvkhfRKLEqJHw8eSk7k3Rh
cx/JSz1t44LOLe5yDA43VMLIJzicFZuYY01+ZMk4DAu6FhIb16xl6oBOShhP7viXrJcsn2kh1Gnj
XUMx8q6lbg2yYw/MF/6dyurGzpANvkYHwaeyQEhhL7G4pfbXypt3hC4QtoQRqUn2rltjxJNs91JB
hsxRaDQ17OVr0KJGB+IX8XFUOpZoG1MCvWmQTjyaq/7rxFEn2yzQ8PKO6iY68CoLKKwHYYRtcIJz
xOEL9A0yknF3AC0+08xRB7iOjmwIVyCzMfDUv6Z5SirWOpv+XCgAPe6HgtjVAaSPRbzrRD428bm4
1JQ1zzVVvqtDGx1es2u4wxW8sY+TDGuLDTzZrD4j5LcEoRl7PuScnj+roy4i/HBUwCJdFB9xqc2a
yvFEzAxgi3Ih43tKdQ72eveLYeC85PTO052GgUN/eGpjgvkmqRW/wDMx7uQsGXf39Rx3zN6nIrp5
bnM9+6/YgHbNPRY7/9Ok6wYtBdh4gJYLmn4UJz9bDmiQV9SPt4TyPEolk/sPCEp9Du8Kif5Ofsoi
V+5xONXhHFAk3UV80g7iPGRQHlohmV37mrZeIdGnrUfFfBiIAXttHGI7zLeW33MQoD4qMnuzoaOZ
njOSi/rz4fIHJetywm75Bn0a546PppDUKuOm17EwYy1b/KADW/HsaoL3kDS33l6fGeWf79WpOpzK
AKAQxQ/SZFBWd1X4AQZ+++8IKbTTsS5YuKlh0lWPlZxMzOHl1VdFhBvLTkzzpGj3JS7ZQj4gmOoy
69VZh9eN8Nco+MHF1KihLkM9dKzDEZxAj7iBEGvtlbQkpxO4R2D76uHc8GDCIU3aGIQFqN1ejoiu
io/Sx6le/MovWjTuA25UK1e1XZElitw7MXe9hdmWNHCbgV9NxeTdRX5VRmdwZpPZ7geywLKTJYWN
vIp2m5/2IznixZuK2eU1oGAshN/noiQ0DRNmbqUOud0oCJFIEh5ZEjWgruX27Nnj3raGE1EC56LD
L/lj9B/gHOz+xGZeuSeJfuI7yCakM0m4/yluSD8aHoWp+TglPwuX0bU4uW4SE+q/DYu9q4uOQke+
FNv8r/5UdUfIB1igb6O12L6slhmL4XN29iDSizQE3tlCrgeABTTzYAQ9mhRZscE3q+qqW+8iwJrT
vm8NBATG6zhsFfe8Uos32GzYKsQy4et63VgGtGlRNmZ1EIcDsocVgNqkAVWdwpns3q9aobbWMFdu
lkJhEYXmQwS5l3MdAKIfGEF/snND02bzrcEBbOJPB3MePQdHYuHeeWObLgRUCCjGKDyXPh0dlzYP
vdC+jGHNCZnGznPTMNJTiGdOqGkoC2H5nptzM4248kPcy24s6s5b/F6xtuFQxMd6Hyh52ygp3Jen
BtLk6tkSfAOHHzswHCbwulFwfWOuqTu3Z+CnumsQdcqYM0OrSSuTWqg7bTwV4nOIjmvpUnYXps+A
uWlSghz9ZUezMExTO4MCGXW5ip0Pjn1UXabG55CdbE3wFSd49cl+GbimY8vR1LY5goCFWQR99xI6
3fHMMQWAIyGhx6/BY4EJDDal+NO/10qIyvUpHfn5upZGkroLnhqcvtfVUwve4Cd/+957cvdvq7Mw
hej9J3OBrS/UYejDQmwyepBPe79cmpf9wHljYT4fzUfBNbm5asz95ufGgJMm05/q8TjSj3b5QMqd
40kZkzuhwQ2IvH8LmxmRYTcXqxeUeyOSguYtMqoqZBvJw1nj9EwsahrUeu8gcot56Y6IIvVd82fS
EQyHtO3vYt1CzWTuoAmomN8KXMSGFWBzueSx+oUqACsej0bW2k6t3FADcnUBpRwkMGQNNcw+K/6k
5nNhfT/gLQFmAP3KdEvljDAdsItR/lUIixxO1twR0s6IdllcJVyWJ+4l393RpHXxKaQe6VPoZAIB
Rbw1Dzq66dnP0vcrC9e2k9JOw47cDW6ship9KVDMVzFlxcIegXC/Vj1LPJRA+iXV4++OzVYUYkoS
qI8vSLlyEGJ3wkfaQ9MuTaH0EbAZxhcgsJsu3MCS+bd8v0LmD4IweErTMlxkl8BCEokCuybpLbY2
xxV6i+8Fiuo4IoncgxbUR/2XZuKQCBLXMywb1nZwvdS6lXQ9i4w6zukIZsH70FlsqE1OTZGuaSDc
XP3iyKG2+qQico4pKz2oTMcSBoEqUeTG95igJUB/K/gwRHrgFfSlB0w9mTkQRdiNnJLNhIc+KXcq
VV370IfLpk65uSnj++b3DRP3ioKNQiahkmiXo+MhHO9V9eeoDQAPH0wx1kY0MlFdhyV3D5vEwQnX
cTjpNG8Ti9XN8DUCd1hBuv7rP7YWoBx/8b/zdmouoFzpfxZ1LlnNG985x0jfmnh066OV7SGBgzPi
exc5JNs6puCILEDp/Bar/3kpulU84si+YUs45o6R3HQBtz5fwlS8NlkDR98g7/C64a3GtpTzQQ+R
/CrhjvUsyfkmz2/axp/w2OpsGMPDkonpKTvM6Q3lxr4XvjQOyffQjHKp8YGWedPKJ9qoeCSntlWw
5+wHxhORVcumoH8P4sBN3YMwzJy7BAb6CHcINktlANfaDmvbMdzYhg26L8Yn1MorJhNBIZc3OYk9
Hiqj9RAqyTkJqwgvMPiUbva7N7+0EpCLGdnpsdia+CWQBo9LsCwW0LTvxeu/IFUKgUO1o147QIso
3MMRKQ6tqvbV7rftoXo1Ex/zzWMTdPj9+rFevlyhYnx+GcTj2Xyaak6JkL6RTOmoVWPJVljRkTY9
9beXQ8oKQgoZjF165L+WjavOVOLTKnsjVin9TSXVNXsw/m7YHrUbUGSiqsHr7UJViBNM978Qno3P
WV7rwzzJfDS3IgCu5EgAxGNh0j1D4h4x1zR21nMYCTJI4cGSIKcknC4BVi7hBGBMKM86X/jeJEqJ
tdgW4csv3Fqk9lp2VSApOpmiApBLr0PXbScv8ihN+azZgVL2u9FGmVX8O/nnHKB6ZGYmaprR0eZ3
Q4kjHBMxEoUuta2GKz6krbB/mFmnrAKhmITXmHwAfpurrhCvcB3hINNXGI/Y6lIZAZGT5qaJdlSR
wB3zazxeKZKJ96hceEB3CH+QX7VuZqIOnVPuIQzCbvZqEanqJPNr0DGOnEAlxkhP72FnqW1nPzhm
iczFEC5wkDMyfBketpDZpRTjlNH1vfpaRQ37L8CHg2LSObpkjNECykQSx4CLP+Kfgq6NcFpy08Lh
+rYLoFXFMrZ+3EH8t8Xm2wOeYRZQhka7eXV8Qrcaq9HSIyezMVVuYiibVROWZOJ7Za4O5fcjLiqh
pX+p0bkPuxlBKxBTAxplO45BHwUp1tCznogY0k5nriYR7JOVBtALFtwvJeGPfsRn3f/n119cAt0J
TpFMv4EVYg28Aduz2G6SCYPcBLBUJGhOwas8NeCGfRCzihirQbnyT9nELmt/DKtv/+AO7THimTiD
mSHVilUIrmJtkhKInVVGjX9i3IqXjIEHYf1fZMfm300CA8TlkYlmy3otWIIG4NBrFGeERAVL+OfF
W2Sy0NMqHnWNu0BYp6MZ4dZCsEWm5of0Gqm5coIMGpYKAIANOykBIUpxCrKGpNQ3FMbGJG3e8kNw
AJVF23j2w1ZH6ei7+zD8OfxWGl0Xzep1wmiYKrWq+6+nzgL3d9sCtRX4SjzXIGtNk4qBE8JV2wNh
yBqObqs1TIHRJHNri7BNRy4CZ302Ziz2cQStB7rpS/tF83cJAODN2wpbe26LH2gqtNsqJzlWUdWK
1JbenVvTv+oitM6RvJUnXw2rKtrd6aZim3V+bO5UeWGhRcKW6K9ej7LjRM3bxRQ4CfR1eEaSJimN
g4/hV3W0tEqsHNou4ckvu+UoyILRhj+Yeg+BYR4btCZU7NNuzSIjgZhjoqNqouGzq+aTqSGq9WRN
2APhfIdHjCVUNFuDm15KMfCasI0yl0mXBkXxv+tZUvZnmYOnGLTgfTWCErThxWvqvXV48oE0YbS2
pMkOFNIUdEQq/pNVzoNPJV8KC8FAUgn1EGabbXR87w2FtYYyndnVcJXPhcScxQoMzXpJLD4+Appy
DCiC1Z1nQBA3Z+XdWfyqAhrBLl5tiEOSRy6GrchOQOyLQcAOiuKXWQ/Q4J2439YfcJTe1yHf7UHj
jTqYRXENJrCdkrlNOGC0KvfMOrDVKMzw+kFo/48Rth33wzC5qFD7odQnYYKFPOEYuiWTrlj/GtRL
mgtedW0ViaZQ1O4vThopd4JvCY2v40DuKSp6wz2yTj2DoittOGjGmbjUkQVkEZ92Q3ANuYB3QKua
6iyG9SsApdEbCOXT1DrHUdvS77u2p4b+rw6UnlFgk8PejKVNMIerxhJa+Jg028NxeD+aBU8H0i8Q
A9KM/eT5R8w0AhXiv73WK7MwvyqNf2HEVrUUVcKHjzBYFeIfXBsybepHx1RX/7YcYaybh+m5POb3
KWSnxZFMkdJZ2HAb9RZjmkKFeOh720Cp6VM1p2e7St4rglOi7/4mAYZfpsLeXJ40++FjNMZRtJk+
RFXYLAFzw+EZi5jP4JIHjdtZvkQF8IRahgi6KpVYec8Iie/NahtSfPcxH01hiUGYgmvgbXf27RRm
JT3VWxyaxFBo3IOZaf6l1Hlj5mZZF3LSCTMKijRxMcHvyda/W2hirFMYuGriEwwkvx3K/pX5Uhlp
1F71L1yqqnbY3wmGdRFS+WKsQ/2Shtp2n76kS3yiBZ4KTjRvGqEIE66rhC5T8F6ucx597cvy8hqj
nVm5DxxHvkL7P+xbwQys1Gd5+3Uxu7bVvftnuM5raKdkYXy4+GGO0/tW2N5X2ymC2NcGbpJeHAc3
WYErjtVEU/J/jxlWLntTzbXnM+AK3sBu3x5cUQUUsOXoffsqxTk5lCfZTRFL7wpxBGx/izmvJ1TV
2jriGX8ozooitxvcPuleAb9dd3uC44gD/BMcRkAxqwLoNDx3viU1r5kRkEoWpg88vBd6gfaRIK5z
npr8uNvBfGSRsB7It/KSqJ32fgHAC2Zg5T3Maa9nt0zz2MCOoL6BSkjyCXEgrrRk3tnFPrKtWoiE
Ji6qObpVxsSUFtQpu9YlaS+7RKfNFUe3vEn3RN1ehwaK8lxh6H54EtNqwyuD3hqkBEWEsYr2oTsH
iGR8250gpTNAwm8fii8ptZuxYvvuxXwzR05IJ/6mwLIeV9lo7uTntyLLgXXBG7aVnwaoAsuGwz/0
ntJujScv07S4Q3aDrnZ0eKThBIrlQspeSE1PwJDiqJbwIlO5UGdYNfc43ikDwt1zPhyrlsHlj4X/
P6hSmmJfimp0tjvB5LSCYJFZgVolJKhoNZ1TByyiy83ZP+fX2NCK8M2HgBdnR/O+TTfhn04ugzuS
MJYfXggFltS0CUtE/wlpIpWn7W9kF4MOcIAuIO+B1mUuh1vF3gvLBf+ybOCYSHNWvj3cjzxa8vHA
qsINpmP/VkDfSc6msj+oJNEULNb+R+qJs4nK8iV9dy+OIPy7jWx+tZoiIBBVFXfGhu0jpJq4Ozob
G0Gmoo4+EFMO4jj0ZtVnE9TbkbcEQrN3a/pS3f3h/IPGn0FCXTFeypxRsoOVfxv4cPRfDbTEl3FQ
UDfHeVYKIwNe7rck6e4awlow2OB3g4RDpN2gvS9UOARz+I1Qiq7uVElqGD1zx5GJulgfCrFY6ShM
najsNlnnyvsLaTBoL+20tXx2FLLTIgSAFAagi2kSuc1F4Tl6VLsb2oEFIgEg0taVd9Jyzx9ogVy+
hEkhbz3f/Yqk5jcDVDsaWQqySvaq058coERzeEdj6tE60CyY7PZcTsq3ZIqswgtxufuqf658xwOn
sSD1vxz8UQW4pA+jCJzgCNAIE/qKTP83T0nlj49TTatlux6b14kpOns+ApOsm+dNgPggQkhBPTUR
oqkr/wMaKa2V/TuwRtRx8NwkuB4TIczLQVq5NJQ8VKXipfQzrFJhR5jYIYjHSW9e0yoW1jlcXDjY
40m9W/MYLNdqrsFSzvXNvEAi3JHSrv60KjWwNCuUiL1wETHKMMVuG4ge/8HhFq/aC3lQ4U/bSQvh
nXzxhIggyg1lRZOnCl/ChrxYJSyku32aGRY0h0GZIQb+D0tb6IpF8Bdi7Gv7lJ1CLsfk7JVhFM96
c6bXfjWDtxtXfBa82rf8x3bxQDpRtoruuGhCR/6l57rBTSn17jl6svkajvaOdpIDot1SzvdEjbyW
07ZlZbbO0iPRxzK2/BSAW2/fahRt/R8wkrkFwFeJxMpeVdkusi5Fbz0+gBMLnSxm9a0GMtzHcQRZ
0nCuLnL7Mmj8JAhAHtc5pFrzOtcLKzh/s81vOeSNaxpJYULCjobApvwu3vuuY5HUo9MTNZVedLJr
seBaPlVje60Fr/cgSod/UTbfgDXcL7L5dvxXS70Qgjx5wUNbl4e1kdvy6tFflm3YpTGFPtWOV9H6
Sb1TZ6YnvlHwxbe8sErSrH/1otR1PiUfT5aAQIUqV/K5ZQJab+2SvMugdq+7QzOxgdNhoYCJ57mi
FwxOkepl0P5uo+AmCdGfjnaufI2OynXSlt//Gsj8wLWZOnadu1yl6nRd6JWYpGlczlsyz2NQsTJh
61l4ojTdOI4RbwLRY7Rw5+CkSs7ZRPH3l0SmIUWSfNKbcKFIZnaNY1lqV7D2Ku0WG0bwNSLhIuel
P7uhI4ouHOQ2lkdligUgwN/XTWmn6wfWEHaqA+SRrqIPdeXPTJBYe4fE2w1xnxUibAkpE+opoHzr
LJKea4heMdwmH15RT7oAvdN2OQnjjRyyuV1U/NN4G5Qaf5CoXYXgesZFRpBFRqoWxPozNJn95smM
giRlkHy6oSiaRw01nvHl35oJZC0fxkysoRCiOudqdONbiyrEtWwb+kk7RWdCmGZskArAtiQlQshL
CMqjkbvXj6FBRTVhAlTHZNC1x0nKNl04o/w2rvc+h2NecuQoPd7aFjqTRrmVCgWVs40omTyEvl8G
wzLKbbsf+IJgB+gSEHXaUdAyQ2Ibwr+XGOr2CJpn4O40A//vFSTg7asw1Vk8Kj9as+TaUGZuIimd
3gTsynsZ9eamgdtcWkgsnqtdTfdtfQbN7hazONaL3GgzhpnO/z0lW879amoF9ZRnrcwy61hOTAXI
J3woAm4MiL+8YIllJno9QBYlvvh1N5webU5WyoHl53XiZj/lps6JL6AOdKL8zEq/aY8JGuYXaaJq
5mSGBN9+LLb9t2PAOkAIuivakZ0G++iCZSak7aX8kwxqLxtur5VGfCsIlt4JksUV/8OXE4A7oOOF
/ovdvfjyAHdgOxdoT/2RfnDm22+gP1quzeak08bBIs4=
`protect end_protected
