-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
mJPQTxiUHwJh4/R3n0Di951llyntfzSK/QlehJy+1dDr9Kvglr9C0K/gBiiVHOLZNj7TUznWdwzC
9f8m472NcH8IjGwNgyRwb4es1icUjevziAIHVO02635M73WiOblk4cH6WJsKmO97RpiqKWUit7P7
huDhYc5fKsqoASCSoZ+smGDCy2IXZWg2DTOD2Msku0f8ucSq0XpSmmwn9hxRjYz7B2vq0HobXYFp
yBxz5D/dWOi+sLZCO0+ET04fmBKzwOu3XGKC7IERce687FtfiyqdB+uui8//7H5zqmtpSWclPbZR
3HJl6x4HKDXmk5Cv8yly/Wmn0QUJ4SCJRiqXDw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 34832)
`protect data_block
uPGzU4yU17Pbs70N3rn2ZzZwbwgZ2zPDV/75whryV//2GIM+5b2L3f0rVANmedgbQqM9AObbxyBd
ywWC0fI9bGe/GjVDHEfwvBwt/Zdn3fcwgW7UsR8UmbH6Jc1HWDbod0eowXJBXspLJPlBHoCVJF8w
9nNK4d1rRlACFnqe5cBY4wQBU9FWG3QzxJzZk2doEFltaJ0+cWxoGnslc5T0nWICyFytoFCrPlDI
TlzGv5Ew7sM/n0q/kdiAdV3snD4aRbUfKkJN5NWc/WeJ3qnanMWJ0VYvjgxBD2f8Cyay3pWBqRwl
wk2v3N3M0EJzeZG7s5usOS3b3KVmT0plBm9rVKm8TTvvy7HD8362trVebD+dnwAbKu/Ku54+0rqO
Ef2ibOlc2OM/RX8clw0nC9botqINH1gIqHPeJBaeSUOK24eMy8kFSVa60caB+X+T0HrRCaninLGr
n/TaTXADb0uSDCB9qZF/vkyVOH8LvjWyFAUw0UhHYf2C1jVYJiHEoGnkcZzP4fxG4zzHX74e6w1y
rHLnVwALkJH57fT9trP2Vh98ghbaKVsg+LPo8wa7KvLsHIBaH4Bn9nQKGw+haciOxZCLtjZAvjYJ
rHlmsymbolQNPz0DeH/W150VsDGt5agzcGxKb9oY9hQ0ZTy131/RMVVWZ1PoA84rrOUA1SyM8uh3
qaj2GHm4dTNTK2uNIH12+vPTaxOcqG4VvTrOt6gd+cAOIdxv8FTsSWbLP0JaPMzMb1jHX3J1Hd+C
+MIR/F/JzeQv2oXNLpopNbxzgwiNQbEDDk5cLG/BiAgaQqgzYkaA0SSymbEmax9eiVfFEN7g+OU5
UpOQzVV2YQvIyRH4apwZ33NyRIxcc4qZyb6X+cTiaJHpT5PfitE1a038QA0qu5FARzX1yYWAMBAn
K884q6jPBSlvJaU120LboFaULI8HCWC5M87pmYoljJ/14JZmQ1Htr1MIk3RPHktS6RWbZ3Bk1n4R
jMeJl6UB2CflmyPIjB4TCZLHh6z9jbzwD9LN9L+nIqRt/URjdheSdGMJV14NxEIaRcn5ymclxvou
A9xKjckb086L9Gs04sHTnOP9Fju6UcLrYNOYPilf4sL+i8hrfXidxOnqnjfViRJLs2k/Enokvwfa
ubIBkQemuu/Svnpaki93Vj6YGA5iR7Yigy89i9ywiQKgfqwYG9Fxlo1eEDubVLIIW5NF84W9rgEL
UBei9BTvxZLw3qmkDABpLZXBBP2usZGYFSNzxORIU0megQ1jR6URXXtyiGUtoyKRKOy4n2DJbxC5
XArYdJoA5ZhN1AxElRSsFQRhr2DUVP3VkWOLXtWK9hDHFJDgoLk4tHeRO3j36xDVPASIFpJkBHyX
nWdEKvVQfIhUgMYuXw69v7grLQN8qcDMAuavbdXvHcJyNcfwiybwSUFPYSO1HDnrkSuojK+D9N18
SXolZWEaOycd2sJhKSpHjXpXMyRAJZu8C1QEIBtYWFRD0aGvMSoL2KuKgVeLd6WqrJpUGkTi21hG
QR3YNM0/5o0E/yGZy8hDtSb+LlcUAeDTqpjgCNmKT/A6hdXTMmPiOhThG3EHvFnwhb3QixxBqH7X
GEroswM6YRwiwi25v9BDngNzjjzVRQWLogRkoHrHX7Bo4d8ZkFiWy74LFoN8FppS0v4FtppnrTyB
MkVTvhYBbQyS1p1jrRpdDsP03eIT45yU93WsK1MHQtCoHclaxQOaBJqpvbZdoxnnY0HjPC7+Y6As
lH7BVjQsvd0lDMbAd9z4PdoXkloxFwCfrxbGGkCeroKQ1Y2IoGeusKftP7ZjMukKISPs1rIbh7oG
8zE2be/DfFkY9M97Rg7C/yjEIqz2H3h6zHGKl+JZCzHvqH/8mc2244dXg10VbLsnIVSUGYjeA/1n
8Vhn5ORAqdCmC1C/saasSp825kueyx60vjiYvmSY4qqkJgJLQJcUMvaZw/isz/dq401ngNh8R9/C
IHZ4sAV1obxGSE0DHSHpdvUTy14YPWbYdYUBLapNCMLq2U477uYEOPWQ3PFAJX/NE4r/eFB8+Yqq
1irVDh/5oUs3/TK+ePC0757rG35p3yYIc2X/MzzKpq6VKHXfkBvx1a+JXNMo+Jx2WJ7k/FIXCsLW
yHj2jty+GapA3j9Sdt2HJIywCKA0v+Ka1sBir0VYcj0vDGAafeGA8JpaP22LhKuqoM9Yjuu5SunY
vppDGTSOwAoy7wJe6MPHdYMidAb6XWcsyNRdacLY3wtqGAl0S7oTLaeO7tf6O7X1+gGZT7++H1HJ
GGJwhrf2TM8L5DsWpc0J+WXvjcsY/wxnJc7G/p6DhSpGndV6kgvz2utlhbV22bRu9n4P5kWqsstc
oca7l0+4PJr2123UsIc549aRgHgNJz+cCBZ69jkTT9RCz4TaI6w7cv/uruml6aaGZJ+9RnunjJqi
RWFvFu1CtG1GZBs35jMCGzEuIFrVkNxdqSwqWPO6/d/dPRoD1re+y8pQH95qENq+HyFWM+AW37du
+fH98w58yNfN5H6vtogTxlEuFTcGWkdtLLWtEtyEDn4pAIFmq0BbN1suZXjG4rQi4d6rDdR/oVRM
QS3CK/OILnFId9ceVD9t8GWVRy6Lbe7Jsdu5hGIgjm0Vo5Y1isPMrJ6PmhGAHh4fFptZgUQHN7/a
Ayh7/90d58z/ZMk4zSmKrtU1dteKxyAf6/ieXfQ9YZWQRluU2z7+5CbH+MVGVeIdTaS73y8jU8nL
ByP1fT0VBf5jYVmSyDtKMjFSKVwFYzn6MMGLX9PnIehq+k+lyoLvvOw3zpTJWJSl3V7sABDhGR46
5GjnhKVnDupbMUgNVFu0xYBjBSK5Tzt0GQbxq+OBPtoBWE5750uvP/qzbDP9eOg6ELjypFcFet8X
jkdqENGO4Mge0drTIPxsKpVDhAatVm0INjwo18XG4/83pRrp6MgvKaY9UwlVVGEwJTrsAOfSkJAy
X9kPrI25Sozua3knP29b0r9GEX8vLNGfvZ4cxB2u7mAqmISfj/QCcwL6fxV82mnwzQdiWbF4gKtn
D7+RCo4CJ3aN6t8J+L7N2M5FE83VLuyugNblTo3b2C9YprRpQeJcMcROzcgjT/plAFs0qyj46rOm
tU/J5mp0TyJp9s7OA5N9flubEO7+K9tXvyGi0cfO3wRh8UVYuyrbp9eSCtANrTdLpme+K+W2OixM
NcagCi+GGyWOT19VeO7hpeqKDjifxqjJKeGOvqNjdSi0w5Ynl2NEUo2iX57Mzj9unQa26MrDU8vM
6KzWvXzlTMyCU5h1BYYopzXu07yBE/H0lKVuUpGekapNbiVXPmJ0+q0xSIkhwSUWOg9Ieq91mT/t
Enx0uRdZAcbzxh20kylof8cX3fNb2+B7Gl70gYCM2waUGEZnm7zEpvQhav2QCXYU0hQv/dlj2oRO
dRiFO3ZD94GunOGHcihoBwwPYSYR7kQ0BuXwT6dX9Cuo0gOif+9yQAIvy3hD9tlMZCAP05MeJoCj
SliiOak4SfQpt7QRWHBgGVPycgB1p+rdfmRlqjz9KI/Fhob/t/6rSZoBOWDZhLeudfYsGpxNeHVZ
MtPhhCdpLTKcWzcD9Ug1xokpuN5COta2UAWit7UsoCqr9p5Iy/ox4BG4E8QpuMR/RTaipTgV9nrW
nPesV/0qgy+hlp34FIePz8v6x3ybKOhmEpHaRcCW8P8l3IepWyR1XhtEI/3QEW1IKNJkRbEPpOLn
9JSX0jJNhP2bOvqW72d0SkmJOmyqGEp6ipNK1FojEz7vfTirlk7uVwqB/OUwIaiFASdAuqUwmMmL
EHBfOcdNIhTtPlhSz1Ml+3CHOKtJx831Tx7EKiQ+k3UqszRiP0gPz9ic80/IrS9weTJxE58ckkbb
xkp9xu7I1HiNhLScRyy10ISibeqgrn81IQ1LM9i+u5WTkhbszE9OQ7zaNr5EMmrgJhYktwYCbFHC
98IxpkPj5r3q74fHNKi5ZwMQBNbHbnC0NPK6K6QQ6y3pH3bcvuVTot+etHR9I22fxIJUYf3PNm/9
jhFdonbOArvpWvm+m0nCAOhhvQiV+MQ0I0ICv7fDXAWC4YQ8+gHpvHxd1MM9xVXyVkTwvumlO51O
V3S5oX96kiJc8Elg3OV5UwO+qSbSP3Cp+kInuXvg8ap1cVDyllcJOkeGlxx8aZ+0lOSeZqhrVg2j
ZJmObprf1/N8ojmS3aty5+zfDJTtGXVqHM53fGy/4rWP4tBfRXJxBVlS2uDtlHAyZRUzjJx9CrDa
T+uYznd5OTLi985GXnv8Ju4+al4ISkP2bBGynMFFH6/XEZccD3CldzsgmQE69dgqFCVZm0gDeiI5
mRi/miCfCgsKnr0QjcNNyUsO+02XOREiuWyzhrz84b8/fpFArUJL50kGaTMa5Ezyh0Jk3mAFS8Or
ldwsYo8ic1B/fh3eUABEHpNNAJFJnF9f5Qz416qUJi60ZrlYZdlNJhvEAve2IipFzNYH2f/7lnR0
1wlXf2Vy2QHCFI6K+GZavcg6qdIADIdERtNzEhr+86RUSE96Tc3ons+pIe9i9lJem88sw6tMtcQc
zXuei8KbTo0VUVs1FA2A/iIfEe0NXTy5AY5rjlzvEbF5A+H0ID3y//gN1jqm+CES5fJEAwNdyJTO
O91nm59IdcrHTYzwNAIO7ul90OLpidoiiF5D36BAmrdFEzM5AcIYL25CzRF2u7b+5p12wTmzsQM2
6DDlOXeY9rkqM/nSTIW0onU9NqEV0MjsJem3rxKby58Yu9MQLJyJ41PT6aCRGcCN0GpGuRp40L7l
tAU/805hKtxC0M69QmVygYBox1dlUJkIEFe0OTFH7WNWDl59GD6peWs39lQ0wTN9OaZYACjfVUpS
/bA0JbRz61SnT33s7qtgdUNX1lJVWKf/t5w0KMctMJy/kSZLxak4kcW0iEFPIDHWn7yp3n/pM95y
HZasS8esUzkwO295wiMJZxAjN12yE0invpufJgCNOi+KYaiWRzCKM16s8efSXggtwBRFoPu9Spwm
j/Tl0sTxrKQXvWhH1CNrRf1+jNLfQjfZ42HGwDNwHnl/bMfWzb4uoxcIk+k7bhnimtt2Ho9sWUE7
DdtvUHHxHb+1p/WVLkn4Tep/SjzRM4jnP7PDpXMJbVYWV+0mHKYHDX9+31x/tBkkXb3m6fdI/uuK
idWksiClf++7DnhVl/gmg59bmjA+I5/CaWiYbSfraLRUJ/t1ypAXUynfLJdo4vjqnXvxfvxzmhaX
Sfmj06mCvsQG4Br6O0erITdUm39qz2AbkYuegkO0xFkhVDgeDpmyK4bPygADcQ2LnBVuDHDF0ClH
toYZEXfVBXiZomjo8MoADGG//TDcJkQoifwNvq5Y2S4Xxwzl1w2Gqwf/3UlW6m9jL41OaMjWePCD
pQBVeJkVDJEBHOEaGIjMGAZIYxYlZMS+YOkx2AYVcoKOmLzHRThQ5QuPBAe5jPPxr1o0lATIm1dK
Nd271Y0QXx1mR/dAncWMVZdjtGsBq2xkAvlkw060tVWFmQt9B/C4zE1OBJvWAVr8vi7BJIqCYGGw
IMD8VlhWZMKCY3A7d+WrME4wCSL4hBbLSA9Zu8nQBRYNIBNrzsGl8T21sM3DXEgWd5WyaKzBFItz
oRBsPgWp553pu0Ss7T74wZCB8GzAjekijIxuYKsNquo5tRVB07m36JsXotI8rHg4RyoHXQ7ZQogG
+I2SfRG7EMp4cZ8dkEGhjGUdQfPUP0tDSPEEfNRiJPu53sP8vNHNf0P70p0qLPYOx8sDjSGJFMqx
tWayhfZUkEqG7T3jOHgBUtjAE7KOsmme2HflcMkNP/dJzQjudP0yw97AhwO3Obo4XEGZ9XJmaOjC
iB5ZyFKt7iaiB/ESXgdgYqiT+OIMcDz/GSC5ua2hHpGdVH47P7BaADNvVbWx9LF1yfK9/IQpXjlp
9Hd9Xjo6n42tVEDM/vWdNWkXIqlFD5i/HTUtvkVSiXR1cxk6Mtc/LUiZ20v/nyqTS3WFKZ8smB33
V0S9oXF9Af3RGmgQNl5vE8xAysu0GtHiyBTX1EddIQHiK4tz0ANyUG5faTtrcP9V8mrvhd/BeBvP
gOMGLAKR2f7OIrb1CABzMeP7ywsJEgRCKIUhqYV4dLszUFUwHmX+CzH3DVcllD+/iHlgePZvSLte
vDH9QHucWrhw1qne1m0kyUYQpFVU96XP8+0p+phoWyF/xE9scCx+ta/Yk8G2VzcVyy8DxqFTzgPt
PY9BNTVC2QuOOckeHZ35NzBqotf8n2Ox8ymd4HI3RMB5WQ8+a9yL/PtUyb4DG6jgzt9kwFM02xg0
y8aVxHFuihcqkiuLH1nZUdPSmqxuE8OhgI9iPBAnqN73S9Alvpluv3MBIE8n71N3fH2B2NOji1Oz
V5gtc+uO7y2U5OS9dMxVPz/3QDQayJHN2reFNCvjO3lhpr3dqmyf3aQMyZZoXv31wQ7NFUl5pBIr
8n6sI/mxfh26KPe9BSywU1VW+sXCg0TnPm8JxMORPIaH1i05iG10oqNcxFX1Kfa8Mfi4WHZ4DtQ8
A+ZHk2TaMuaLsMPNeZ6tnW9H8bETy62huWXGenmMsb74eu2tS/xz1s9TkaWAsHEMB0v0TYhXdeNn
N8OZ/NAeoIcGKtlDLqMm9zf89AwXDdP5oH0a8E+G1baJQ6TK8md5jaPKJANNGjh3/UZymJpZBk6h
xt7Ll6rIJBRC6QH1gs9NvMee+taPr+CLrQ0bKvLNRxaEtBkHkRtHAaFCHDP4LUX+Q5U+2a0tpxnT
04K0TCjC33myT3M0vp2BoP/mE88MHCmYpsCwcAECBTZQtkpSL21p5ZaOX+bAB/mIOGLooseif8zv
aRwOJLghl6Z7i7CqHSj7PACIShWwtCCKzR7H4PXqBY1rltie74BJPIgwn10wBDnR8mr3gmfCaQ18
hiki6WVnt03Y/KnC2cu1R4Fy2TDcblnN5SBBPbuYlo6FKYurx2Y/Znnd1PB1oqKoWj/Xl2+UffOE
KRiERI1vAzmoUtlEOUDgKYluX0ojZ4R4BEvsrEJ/wSLXH/xy8v/yE9SnoaEzwti/I9naIscHbgE7
H5djwkqSiO+KcPEjFF04FCrop7KLt/UNBoSSXYm+v0zqtZaobTDFbKqz+qglpvHDQ1MhxcNxX37L
ZvqBp/zfHjlC9myS7YHGu+lpIn/h7pg65m/YBGqTdk5lu6f5Y7sNTJ5KNWz2JgM9LJ6lv2lWUegu
MSNiVFJFbCbO/WGXAL9HGJLzIqDPe3Iy1/q9c09psk1kEGNU6BuxY2dWZVQZIRtLRpcOA6yRowMj
md3kMA0MRzjMjAOZ3jKNR4C+xyyEF3HYR41BgGu/vW/Fb48csBA6sdpDcojGIMXaWBHV70+Rg1oD
w51Acbg7kdNtDpOO2q1at0AP2eTQSWIq76bv+ktXMRavAvyQOxnZ5pifcS4JjBCesxjIfU03UnIN
iJS39ueFE1T6B5ws/rVBbsQVsSH2Ugr7KwF9HFJ3gde4d2A5X8My8T6ODfOYeyLAXlagFX7u8qQG
hQOmCUnOPQVNhmPaR1DCHv+iU9djBEVIHJT8Hh7ovNOuVwH5Z+SjFIVorlAgItQw+Q7risphjxlG
OA7kV5Us3Y2wCb6bE78Q5dRpyFUbDefTCJVKN4RAau+MffeYbabmTBikmXIdfjbIDmBj3IzRkZAs
ZhLrhmBiA3+0hekXb4TGdxSXwbA5rs5iDiqxP4XMzbCxcgBI1WBlRSdCCsViupMd9bHirf182QY6
vFDFe7Y1Do36A8f+yQ5C/ihbWxOAu446GfCjhiV9ZUqEZBWTCevOnVv960X5J0NGakEAfzR+2Bm/
OToejSz8NfnAai9JbY/EaKtEPBkAS4ex6hCyyFKlIDC9qnrfTQChKxhYjdg6oM6PUO3PCdoUAHnD
73JRCs6iRm8J3EmhvENt9q7QGKWp6q7OqOXa0M82ER/9MTTJ3iFjIPQR6m4Ffm7nSAvM51KECOMD
pmDnmwFxH4pfBY43EgGLBgtXarxM693LOzGICcyxhlXJCBXWgc+ahunJU5TJXC4LxzAD6ZG6Zp/L
GGWy6AI8gsM1N7YtpB02bkm0oCJitVg/frN3E5MlOBpeMDYoH5XkAPCyFDksbPoVefvOFj8fDV4C
USWWEcCJ+BUv+iqUt7tSQh1zWNMSHVNO9h0wOslU+ruU8uYfR0p3/QGKKNbwCptJ4fdrONFF/RYV
TSWWJTHeBafY8Ybz+s+vyV3fs5RNObXPSYtSEC2lTWkxwDyPhg7wr3AC36p4/jhFZoyqGH3VDxTr
l5p8kfs8d/Db208FVIC7NVP0aNS7pMQpsiSvbnM0091N4sxGYf3wQAOkn+UhUkPpZRnz0/pCKuFS
iCypY/CUx6pGbttYCAyKLEZNeJOv2GD8+nU3mB2YgyC2u2BmwRNLq2yI8Cqoi5+ueUYfRlLDaGsw
Mxl2DAUfFVDKA/mrdoiRzwDrX5sJfvRihSmoyfQ984tofCJNdgWKKPeABipUoqZODUaNIYhp2a9X
5zMB84wsO+rfqnzw/yY5mEyZJPnPwLE95gCZH5OYrkWgJtAtOYgOBqmIhSLKd7EPFTFkAqj00Sx3
SOVY6kBqguMxB6Knbl8fJU+m2dYPX9zsPxOP8KZmTCHCVYpsFmPl/qj8KA22mrKTNGAgOvbXjJ2a
Vj8SapImBwlX8p9sOWBCghIF/84AWMpcq/rw+NMYPqduGbzM/kevjSBfWm8TA5Snyj8Y9Rcjl9Ek
0GcXFxq/92XBLiyRLRGmUOKWpK0SqbVjNp0uGfKdAG23OFfMyI4WqmLCezbL8yFyo4i3sdta2++d
C9syXej6X3NHsUy0V6C7gSTGGsETKO1fNvv8J5ow4SFPM4cjVlgltaKSTYsBami1eol55tCOH4Fs
eSKdAfphG+8F/VgIQJfFEO1CeR3vxqJcvpbL/6w35pdRX234CWZVL5ApQ/huc27eNkLZBoAFFnP6
jNi5dDgx/PDC+ZdiFI6UEEFZeFxXjmkeiiOOZRX+bOuWq+5mhKdBO0T/khWR6QlfRhKealigNS6p
XP9rjTApJmL97KHrA5A9HTo2BWA5uIMkwnMiEBRp5vKp692/+YKnmPCBxS2F5Uy6tm5v6P1XmQ52
hqqj7swYD5/XhQP6pLTHLQjfjpTDieyGFEDvN+RWZuqg4yorj7ghrUBJU6qAaxxFupN0jlzUQAML
6pNrHTNvA2UXXKE1nrFTevSzFN2k7j5gpjEcc63EGSs4ra4aP06gIDOs2030BwT2Bs9D4+QS7bPm
Q70q6he1FVBMGAtfmKbBwxQBK+9eclFiHuSztrxJDQMscYkiYUzE0FfoXr4Fau7O/2LbdWu1Gk7t
SdR5k7/kewdiNyAipnnyWqUJYqO4IbRxhZWq9qQ4tr6zlYUGXTa0adDwJUN+ylHpvYw425IsTCu9
WSWSQUh0DiEjM5w46hjy0Y5qIWHw1/cRQJSDOLEjjEpVutM2ocOJOcP0bh0YvWWMKrYb6wLgokGx
lPOTliv1vCLDhbbmD/RuaHLEfyg2BltPLeM+t3IlQTqNBXXQfFBwpKQ4iVc2xsTLo1eXMwxXDqcJ
f2tn18BdUej+OjeuhQMzDnPRo1hx3y0cK/fs0ie0e+ChxDp77YoCEDa6sDmiN4EQU3A+IbL2lU19
EaLy4LGjzuZ6dWCm5Kv9c/rTFNC5lWS1RI+izdsHnagyK3HLxfkevbUuIfBEwGAur/bxvaRQmwcK
pqhwO5TqJP/6VtDAyY+pGA5oKMZDURfCi7cmaXD4mqC05K6FViMZGc2muPimWlJGt1jZrUxP6YnY
kzQTkuMdDVeZNgc6FAOOk9AbmuTFzTblmJML8VOKTCVN3Eqeg/fEYO11WvyaDRsHlBnbcwBwS+kH
xbQrAZr8edP1TNbbyVSpQhxKY8TtPtcG9re0CHoek0o5N1mmlG5wWamFWxwLsxdyyTibfYW7f89y
ldih+IdcjyW/xt2vTiIYifcpdurcx789iK8jV98Gpn3TvTar5JVEuWmMoDLHqy4hXq3XcUgOFEix
5jtE/aTPZPHFoNqH5e6m8brpCtPBV1kI/fZAcCuVpCKQZ6zZXVDSLh9XE4BBGmnECr8iSfWvEl2k
q3fgM62C7BrJxO7flH6vJTkY/qo3+zH+IZAgS25NXt9Ng/z/UgMJ5GaioBTkBnjl0x2Dr0qSypsH
+bm3qnv6r2iEFpuuVGLsmVTKcV1097gcuU1Xq1PQMC4oSuwoP+XXvXNz55Eer0f/so2IgdfDFkcg
nReRITWlKM9Uz0S5y7yhVn/Xp8N7l7gx5hZIhUesjaBSjwYBKP70SIqQ6oFIDvcX0PtmW3KHgDDn
PJ6R3xgtzs/kHo3TXH179gpz2sHNJ1qfMxW8KcxSglGfeSlC0xROnDrXDnaRYuxjY63MK5a82Rww
T12E9GmGOnoJle71zlOlnMRdtOpG+SJ4ONqgIAwsASxRkYek482VzCwdrUCsqcw9alPLMS2b2PF8
nNxLDA4BEVHX4Bk4NtfN2ufKUEhMxZnuROzaCmwrdN5ybzjC+IkhNr10PeQq3817+cAwLwEAGqeX
bzk/73sA8a2eiO60eQtU4Ph0rH78d7cEldZ1Qsvs6twj7IsH+Naw6ilEWTtZIYgPwfXVnn+nBQAC
ODpue5POL5SEPIC62QLqZtMFaADgBWqwhqcOBF863vrHfdudwnrs2mE/XiGSAMgjVPpZjRljkRMQ
zaJu7BM7Zad7R0BKRTEyJAXq7ESdjmMFRG1bUmdwvObdNi9JVUuXk5huPYBW0hiLY5eYKMz9B/yo
KrtRAy3txwW+GLAvDSRSTy0gTlC8RETjpYKyLQAF0wEPcoMdeETsxsr7GJxsC1tnUJgEMwivUFn7
RjbOSaWeQ/8PiriUPmpV6L6HER5qNmmUYcFnagFkti/v6FuXFnHWGMUE+dWmMFa0eTa2vi+MqRPS
LB81NbQxgrETYZc5yDcR1j7Pl7hzjIu7LuyfFBXqFZoDEV1I2ZkU5b4m85ZVECMn6Bu+uqk8dtpd
5uB53iQ5M7QeEVhHy3YMBWJoGAr0Dv1Exq7tju+prA0AgRj92sw9EmLDLbLQv//fOucaN5WhHIiZ
PLUtAAaWuMpSVJcIOtiumc2o7VCAjG9/TYMxyB5ekQKVqyBfCE/UKOL0ZT02PAkO9X0XBCfpIRUB
I757IWiqwwVFrc2g01hAbBJ0h0EgXe27ZUxoNF1nLPwU/dF8+m7k7H35wW8CqpDZ1aVmBJxI1rZM
MdK6hAJ6A0eeQRSmzPHUrBqwbrpWqHcgw2OX3hBM1rGkiM0l8iiREKPd3KYlwqMSuRqFokPJ6yzK
gKCc3v3PxQSlsFu9JENzF0csO5QX8zv7Aqb4KF11ukr5RKTBkfMAzhfAMsm/OQpJl4eE5gqKLPTb
6r9guOLrZ3hZwNtloAh+uKHwlsA3MdnTR2Zy01nPDUWcOLxz7Ov9WKWu9uOdcF6a/MvRZeUStw5x
z8rwz9e/igjZ+cGMQyhKkz/rkUcBK3xYRrhN2fds4fFLlIjbM1myIP0u3kQZkiD1FwIoGuftz4vf
0kobr4mWnpOhpvUHFMQDfeaCe4mJeF2OeLjfK8tSIGxQj+42K7OWBArNinx6qhClMv/57MIeORAq
+qL2n/tunM+yPQ7Bs7RTke1f9BgTmL0Ke1Kj9BgHkE0yPEjcyGJfoX3UHDEX/dYlefrGNZGSV31g
C2Ff9JADaLTdlPk+3ecE2+/bxt0Rj8Fa6+WsEHE+1uirCXKEEp3izwUC8cIFKh6u/HV+Y8aJzM1P
/Bt1JrBidRftPAU4nKIwD+HNa8tLrJ6QietYlt253enSDvTwMmtXJN96va1RE71xBjY39/t+GoSk
NGUNfUyLKWruZeKK5rsCMPHXfd/78iyvpleO6ShFXi3McpndbO/3k4Nou8flUM+vRua6UfidDujE
OvJOba/6DpAIss2BziqaJAur1EFYXncPSpHUV1gBXuWp3JEk5iIPp4sge1Epobqh2tS0wYEUQJEr
+VWHTJ3WNrKndSWaugOY7Bk/VK0WTLoDeRbQKGb3wgsXG3fSmRUZSEmmxzzpDhVvSi8EwUqY/sIU
o5Q40gHXHWocksNEYhqK1Suq0NdVmTrPmI216pY2Uc+jnZrVCFw7eLr+QKLyofzr+emTdLrK1QtA
0MHKT/qnJ/k7ABUgYaRliTgQR3phNcuQr9fAwhHn8mibhSPfIWc9cUfliDOEvRPFcJMF8aUgrwak
m9vLfgBGvmoj4UGCElnHWV2B/hS0bkJOSBXii8yApSrItlTHuuTQxkGwLJRUU1VWI5rO5GRC32dS
WKtYpeTd1wfkmMKv7pvEoQlGx4r9AcTF8NP+haFDbbpzOrhSkt6dLK+nZMm0qcruMuEKEpVriozR
1mPGoPqWwc7kQHYZvW2q5yZz7vQBqJPQqXnnhKM6Rr0Hoj5kgvF9jqA8DNyAHb6N7QitI0SLRowG
fAgZjsVjp75Tqb4mGirQPZCrpntCfokedUQa760kVUkqT6OlS4sekYEQKs86V6uqVOIIa/DPzqBL
1HFmVIJKvotLzj66D52HEPnhmdtfcw16XefRAc8qwI/3EITZbmCNe4SOhC2uzLxPa+Dr5a5rcPMd
FJscBSneIRTf0mnu+TbievJ72boMKdNy5LglIaXiUX1KBGkwkqi9CHJaPKjipxSnkI5tQ5FZf8Zk
ZQn/XFjvgpa8wEDODNOlhJpLlo4t90EY3/5fZuc3n7aX++8ZGSX5TNIevEYpRVmyXPnp4ES/JeDi
pOf4dtl2VLep3uczlgDzbihgFsw6KF8zQysGEPtC0FHIH9kqhhtkr5PFGruPVquf5bu88h2cBijj
+5CbglXl+kALl/C+lgOghlN/OxabUBD7aAuQ5QQHCyplPOi2Cdvbwgnu9C/gQMjKjP1bRCuzEKeE
4irLx+vmbJxp3lkg3KnL+gUP79Vj18g5qrxlESh/yY3/o2ER6SSktzaYVrfYQ6jfGPYWX2TRKdbc
xkJIiK4sh4ixU0jqWujknoRXKdXMcTctO8zfVUY7pM4mMf5CbV0y/Mv5772NPqwX4y8CTFZTuC0Y
yvlN8wg0MBYtXkusbZ9kwGdLjw22LENxbILjlXoDUvhNQj9a7okRGpRvIrDIsg0q6n5Rfxjz70j9
P4l4ROsUtiFscFII5NSOOfb9ec4pelSokvso+RTrBcvwgrjUQdll9Aj0zWQJbFk2kPmfgzNzM6w5
5d44Lr01cBySuRUHKkgavdQlYZd7ToyAftG0sPPjRGkzw+xl5qHa0D/2KOs+0ynz4lXjXxCArduj
uZ3tNIhJvFbJyrCxgDIqRSenUunlG0PH7XnhWUpx4C5yTnWRyNTGxlvSWU+wyHb/AWwbnie7sTS5
wcFZCubtgFXORI0505BYE2uEXjabA5YysBq6uiitXvYlcBoBZaBAWKvnP/v+brMgaStSO1op2rr6
jk0mJDaIMCHZH8RgfD0SWDEduecniEt2qtmp0bmx1Im/4z6AfwfH95Sq4lITLm5PCyTegdTmdgwS
ID+hN97sFYPCPynjo5wfzNlGADJSH9cjZDnH6T9REqTK3lYLzMgnF5Ai7GpyHC6gv7538InIgTtC
xOhcHkKEuQD21n865jjeTsGufK1TGGpdhYYKhfCAPjpw2UZW49SMKH/6lAKRLf9yK06flHto7Ud5
vZiMRHRgKj1tNHTdfrQb/IWn3ErCDRcEuD9sB7usaMyLDACLdFY1APOgVq9b5lifFaqRbX+0OU79
juQJamWSYpboKP9eCEQvo9lGgfF1Dkq4o5moKTc+rEXH10yYS1xPtZ3ixPfKRgvwXiuZlnerw0Gh
XIUJUZpyMZrCQ4GIKgU+ldvJB9ZMRWgfxG+f05YpAlwV3KOl4OOmyO3DNwZhmTq/A1al+IC6zltG
2aJJYQ/QzX+n2payfv0TG46ZuSVZ5/2jsVWXF/487FNI/Py2frbU43RfYn+r7hQ0nn0x5uKVbTD0
A+yKlutqUJJGaeAQXk7s+4AlcCZxSfOqNXRvE0Qc9nsie0X/1AKyfFm7JLgDEyH7ddzUBp1/9iNM
F+yjaXyEZkKnTpO+HJLSu/jytdOQNnZcypjgqnUbgNfZ6vD61v4LL1OdvlLFHqhhw6WIgI375N4e
Va+N2fEZTSvC4Hqm4/h3fo2CkvX3QM+aPhXBXy0ROZZPWkL/57+g82nNbegu04E0FuecSjFdvLLt
TmyDZ/pgot4fubfXwSLFHICMRkkbqUk89ybi0QFlEUjUX87Fni4m1cYNiJ95qQlaaA1m8FZFRHYO
UzpwEUaES2vYD3smKm+Y/cxq1T4Mo6zQbzTuZYIJiYHDM41mIN8/93YKnoxrLHPDylByH8J0IAxf
JSh9oIxnpaqB66vYaJQWDE54mpTFeyWoDRj2hZ5ddUnX6J+L6mJ/5fNrCvew/zkbxb70R2MxkYph
0GRPpjUCt8Im+pQS218vEhGbqCQJGA6bEj0/0lBvsqJMI9RaL6SesOIEx67tORINbAYylKjusrTO
YYioXQ2ygfKmytehU2ZZe8Cy9Z4W4PgZxl8UNBfN29HnKb/vmaeaUmqRxhl4+heHSl/rIDmr9PT+
FqnehT3cVtmLxHYEgtZSLIb6f28tXCjAEDguSiunkvrLT4cRLiPSs24V/BgDl/s/7imk3rTm66M8
fuoCIWdkaEpiH0bgSlTCbmD5Yse01uWonpJX0mIrTCyDfBye9GqlE56iCQSRHUiQ79HmEWyN3uvi
BZXG1QKVXNsBShJ2PuOVIJ8DckNED1KpPKswe0yhLT3yDranb2cG9zjckidPkC+VcuzTcvoU6ydn
Dsmp/khv++6ILhiehJYh0lLAahOhL+6dmqlL0RysPhstRpXUXh+43o7Q1gyW/KljUgPQ+L+RfJmb
huFrYhkX4GiOWfOspwngHtnrzYOi1rLItUoSRhgI65hBiuxQZxjlxMyxZqAbVlxOhn4ar35O2i1c
dl/IaBEEFRl/7cxxyfhUQnYjRIUTgSMFuqbij8DtkF68TcZ5+J16Mg2YCZ5RKa0h0j+b4QT6qv5P
PZ0UQdHRMVdX9aa2RIrkGcE0mcpm4ADwbm6V3ViiOxJPhe5P9y5dM9q7SMeUq+97h6f3vr8Re9fr
ncR9YFV/bA9TsUboBH752jP9qoeuKfeHuIpQiuXZXdoipgUTHosCcvPac0RRITXh3AebTdi7at81
aiPhC9wFDGYa8mhyxhJl6TCpTSZP6YidCimxAMLP04ELPCyA6192LNbMyQKTUocFc3zpXa66HsjH
gky6j2rmjC9cZAyYBBaAod5doK/yo7GMHIxPXmoVjilUtgLxV55ZALQYObjcIHQfwpyU92ZLJqNC
diJmklGzEtwCsT5GNTR++DM6seBq8sOudpx4M2EnXHP2Lo9n2pdGct8qxZbUUgHzJEKmq4QgkiDd
XM3vHWOvTWGl1USkj/dhbll2Y4zAb8KNVhJ0y5J/bTMEci8FWLesj6gH5UQcnMwACP9WxvUvS7Ii
wBHKGHdc+H8boOy5K+d/ZqPiQteulVHHsaexBW76P774Y25w0BIBxJuPJ73Oyzg96CAKq4u0/7I+
b+JGUm1NSf+pZHjMOl+HQHBFBzo8F6ZKjAwmCpDSUZXVyXSTVsqLHmFOp8wgnOehKPNo0z4brBrH
sHIxC1DcDA+x3GfQtUjRa1N4ilTMJbmma8Gex3NfDLjPnQKuDm6AkWUkCdHeSNjkwGLeMYk1838+
iX7R4visSzpJe0Uc6vU5PLC/5kr3s6qUXffq7oHuWJ9G/uV9GzEdmkKt5U70/Jybrsh2BcU1fDVX
bxaPstl7HugK0D2EclM2KudmrtjBYV2Xgkr7N5oyAFX0axL7CDCdJlL+6/3ab0ijJy5Y2smlIXCs
OTggTsBLFiLEVd1bpAGxGxBciwY/v7BtUDixWG5rr7bF95c3DBx45hnzoi0sSgWYGZSO//L8UYSm
TNWYIpsD8h84j0bhWNkRyzIEZ5/WYlLmLr5Ewhab1cjDPOQwCJWkSouY9kVRmzy4jD0o90HbVJhi
Qh/972gjUi+vIbhuKxkIU2XUGAOPKqBOAoM6VDYE7KhUzdPGRIrDBRJBj8+4qM5bBtRxSLqIRGw2
My99uzm8MyTM20hznzoDxT+TZzhdtPx05mAeU2tBEFtJYPxoe/4ieIqUG2E91j0FC/HWSrNUbZch
OFdW51WSPmkTTVXXrsOCJuS2R6oqwJ9MnPuf6saia8GBCQumx4DDIDMUHdIDan+B+Rkq+2ArIV/k
hpqOl8lfn4bcsmc4Dg9ujgbQpOxwhpMjgMKKzXdoGL/PUkiWJcvZwmDOfTqHfAZLiGfR4lXzzw69
ByBisRXUyHRwfmVgnPBHzKQqzhE5kiUjCXqCq+T+TpvupVnNDOwzXSf+aVv9B8kfoDtwDhPnO3I7
wC8qbNpMlHlxam/RQ/fDMoh48LmMioSVCvDnLFFeK685YnALRzKim8gMNrn3wsGN5NVOnkTwbpO+
J6wkEFfSsyEpL2fWZvfC9zp1vrJ6E0usZzxeDmOIPrOeJa+iJe98zTX2zFH6+O4WKwFjke/2EdJR
MgteWdfaMiqyk7C3L5FAY8poxHNW2E/KeasVtFIMYaGXix23pNiVsHYRxKDz37PNotQg4DqP1SzU
Y0wkIK1TcdkPOH1HaixhgyQA9+a+S4LYXV6MPPQAo+j34pekpy6zIF1rwPa7anC7HsheSIN0lTU0
15rkZtFl5X/se7Ql2zkNs69j/VVzi5IYPLiatyDlmwb5CTAj2GRwiHO3Wlm5t3OraRoGLE5sPKTB
oM1i0EKRkYBWmT/koqwqNHCWJLZ1O+zqXdlB7VkBtPyoHt3IrnybRUzJDXYpiGq+Gjeh21dOjIQu
BRdvJTsoFHeOoX/Vtfzd85AXwQIghgOcRCbWBBX0/qVligVAgvomKT5B1aOXXB4VvVTlWfONBKL7
pKAzRKqk2K99YzxGcTyYxD2/VhUdgSlNwAYMUXo0MPPBea+vyXpCmvlBmPIZAVJ45f+kAwRFRTkm
IJA+oLKJVj4Dk7rX6mK0KO4QpkPOzkrjG20DT1dWE+JABFxn2PjTGjo3vaKdhAcq9dZKpIgniFeJ
8gU+Z7O5fKuhF7CCd8gZU0sxlc/ZNHdDZJ4P+anQ4CnIeZxVemqqgdnj/0qXSCY7FBwpS+/pHpM5
I/hRvSVtHHr29ApbkvibOVIxWC6XlqHebttNqM0gDjcOl6Fv+KIoCfyqRUbDWdtNyx1G+Cp9jKKY
26tfGyZEGe8ZIZnRlWuZ8r0yt7PN8gaGSi1ACWr+wIEwVf+b9BkijN4lBo5TOhwoowYb9aszKZ3M
l4QclKKzTQ98K1iQAItFHw5jkq5XVrCbZZ/+7gWyTOzbMTrnv1yGT8hPoX0Z6rOlW7ZwFix1Bqnp
tnWUsLziBdAyFq/jkTxciBBZpUwcOL7nuQhDZgI9uWnsdjJaCcY04qtBfKx+8PPEM5SF1bIuzjVM
01BtxKhlh8KFifZyTRy67fJAeuwruXrO2hGUPB8PL4hSOFT0FpjJ5ABTTnJ2tFvVbd3Omz/5mHy3
+PpfdPo3ZxIDlEfZQZorTEisNRRHy/xZsOJ2gxHFkMZpaT9ACCX/pOTmI4huDNDNGdOgVUxuiAxe
aPzNRLyHgcuaUdOjJbkdibYq67luMoJqAUn9ObdargN/sBBCBN6z0G1nNOe2bSb5vzqz7nK49KnQ
1OxdkViPzIqYZFYD4zCIqhelx+9Zi8YkHBZOtOd5vA/GL8FVd3o8DD5+ICSskuM1YLzoVFbFwDNw
mJ++BY9ponGxTlVR8wycTX12PpIuecw/M9gfXEPtH+L0VP19wFgpWbx6BoVpj97coLSkx4UwNrzr
wL1w+SIX85y2tcWQRSYyFsDkbkqt/s6CADQzQ9qx7SfOygItQ/IW3YQoFEjY9lvTiEA8GX1Lus+j
gNC5fcTTmGiFI3523dK6DlR+p8xPqBMh0HWqJQZYDKHXRBbgjTkPmaVU5gVes0SivAaNhuvmZRfn
7B2KhN9sZHGJOIJHaf4oSfD6jEUYM7vlz3Jai5z3axMKR0H+XQwbp3koQoEaeeI4HWf/wnoA2CHE
c5zPanp+TZcuDcThKsPJee++GaqZoRM26XA5Eda/iO4ar/B4D/HbmQzccAm7Ki+fX1S7vGvkLSTw
BLBYrkFh9XrLXkLmGcyocLu1Y4cNzAhrWmMoqDTt+nOmqNLs1qmriaUpiCUvpW/zjy7wSWy1iE9u
PobGIj+XSn6QGVUTZrhmc2q3x9RkNhIrfaub67peIQyYobNx9dsO2CHOLfi2wVjHwZhnOn6OnOTz
vHnRs8SIHvsUyUGJ6NBGl78ZBXl458NBz9Q8K/gCi/U5iNmW+TjSrVtLLl1W69H/3dm2pQaeQyzX
LfhZYJ4ItseJ/oGvXq5mzRSI1rm03tJi/tBEzYstkI3V2rfXX/fTWL+lcZHUdLsHX7IBqFGCplI1
Z+dWf0tPSwWsfri0WeO//27CHzkbgh+IAkj6rtYKXCGimyzPowRMLvyGKWqR/z2bTwvHjmfziD/r
Tp2w6CU3bzNFhM+JeocJzYET8KTzoC+utRF5ph45ix1xfn5Eynm5dKrPh1BhvPRBBSrFBW7O0ry3
tYAMtAnF30NFIawXSVqBC+8NPpWfNnlOHysZ7c48yAUr0+lKwirw6Uv/29YNkupj/JPOmsSAvvvj
6O1JXyHzW8x0u57PZ9PkWi8XJGeoiAcg2OmGJCSvkmhU7QPvJVQ0LqTeeOSnNnRcPyh+fdK7QHH2
kYnftrhlb2cvofoubf2P4197RdVXMUpQ+rfszektBQXC12CpC6wAPNF6gXFlxugA+CMaQrtB0luW
ZaojLgL6OosdT45i+UHSVrcC41pVnnCGljQ5uUklh4UuT/pIChyoZ6JplItqTFR7SIDgx98AmS8R
bebZ8j2uTiXM0pIk5ATkS0u2E9hB4zEn+DzN/oHvt651Yi8JyPKnGh6WyjjnVgZFFi+jyn5u0FQ8
yDpxmEMkq3qrVX4T+1sf85A1+5Cul7QuaoBdZ1DnJ5JnW8J4uv1z2kWR+BPBQIcDtB0qti9VZD7c
TpttVymRNcCfhftAv7WyxC4Wj5ZkZgyC1GNwf6nZtcokI2asKB7EpzEzutphccCnxY5xYHMlunvO
xiVWqhgvnMxismDfKS06kdTESkkrfgIyuKowp8rpfL6Xs3DM+pqO96ycUb53ElpXoU+D5WToYzC8
cYn+VRZu5OXKcs9myhOov+wYwhnaXVfVK5PaW/rnbqJlRhmS4uK+u+yvy+K40WtLmJBx1sWkFrH4
tlSUKAWkWVXFZ15mrxXk+1xFlimGXmvASeGrd0BLgpFEZHcmSBvHfx9nHYzgK/eRji50lR5q+Z0B
pxwFkE6YoKE8lCGYSngCL59LP4FRv+Be4uRf3e2vaibgf82i8vAV/vTRa6ad9mAW5RX1HLGW3cPe
jHv8xR21dDFslit/R4CttJDhOb+6vTJ8uzyXsYBndhmACeioOqXRN4a8ikJf0YRiFDOT6xb/yubk
oQdw4on30kFnK679tEOOF6giDvktL6eWS/StKuzu5xypie6PidPuqU8eGqx879PKBCbTCgaV3KqZ
hxiYN0F/klQkOWP5Kz3jQObJwM6kdAH/weGBCMA5gT5PfRp6f+Dw08GcOGGvUXfsgBfS3Kq9eVbs
B1rM6bTKadyjTQ7shnhn0L1B45cO0MjWNC4CHSh329jlAAqRFJUDFP7rJR6y6M5uBgQnYCuVK1LW
Hp437mOGkiEAfIrgo7/VDOfkwXDnkwkkcD1iI+IMY1L0PN66GegSsd1VH+5ktyj0PHRm5tTp1cUg
Fi2OkBsltaRnIWndzXXjrqzMXki0uzogK2GfyXXsTWrVfy1kQ7Mq7XOY0+g9wUHECP+uxnyAvYNo
PM8+1V1icUbXhooAgoeQZCEDku2xEaZgRmCbQ9X82KPz2f0WwQFZ/vxBJ7aSzzh8l/Jed8Tm81Rx
Rq7yg3fcRBDdwsusZsXJ6E5kt9YUbo+B6FAZIF3EHTeS7j9grszw58OTWQa17EISGceK4nQH9iwY
aihGRHEt1L4W1qkDaGbv9j+lBmB34dOg3+Q2AG2Jat5YhBYd9qHEmyQIgINS99KgZhxucvZM7lKQ
oShVw+HMRekoXDlXdoZHEm5DdRH9HHTpLMScK8u4R7vCkURwumcms0vlf2UPuCNSfGUgFzHiM9pi
MHS7FPsPZrwy0KcfLqnGseT32boin0jxSvYefU3FQQUmQ9oqDYF02foEGM+jxIG5/sKwMFMwYDdb
+nYgHXMAIFWkZE+9fc6h9891JTvSaEjQrGi06WiOBDrT0Zxhz/SsrlmaduRTh2KHCSS4P4Ii2h4k
eyG0UL5VwqG38Mu603fDlVYehDsu8/ePK9A1wjN4xIORagVXnRiUuuf+SqZa7JXMV5HlNxDxt3IC
6iH46R5raOv4T+1nmXPMyK7bZZh+0KTxhntQEAF5lGOIET6npeARzxZ15j1/VKC2yhxo1UwxC7+a
ypOrdEIQuvOuSf984IvRnWHr8nQM44qMgadVIxiQ0cuAG69uNmKrkjmauE/FYWcpuWsgqxaZdZjR
c0HfppVFGqXVe2p+pZGZQHRbBfhewWWFMWFOZDSVuIdtDmV6jIf52Zt2yVk+TSqJ97N+uavRb4Iy
zc8+9Ka0m/F3+7TiFgVD4aSnilE/DvBMCSpX+ktENbUz+VV8sUxLo4goCdn+D196RtrNAnA1Y6Tm
HU96mTrRU7LOu1CgMCYkN5AzPslkhejUo1/QhyC1i+ItsPm15Q7hf4gYjo/Gs+lwCq3eli+sgQxi
PoQPuiOFixKuOS7qtOs1o8ocNvuxTy3XoCk1lLY6LA8bLYYVAJHxKALo72qjHr/vKxkTMQtH44Ma
fnXTrVzf0pCYht1vZdqDyvne7zEXDQbRGPM13FPQ4rrLIHOffsuqiCoCGILNuhKOLOohk0Bq/qcD
RvYlYJ8z4HRqq3Qf4fj4HNmjc318ApENnp2DK5/0/wem8zh38MbhF7/OBmIUQM7VgrESw3iSykVM
oKOmnQ+bZho8fP505h3rnK9tDy7yjwyYhvV4lmYiammWcmLNuL3EmcYo/x5lI2Q8ShE9vmQy4hIn
WuR7po0Z0gK0QMq9pzmYRW5ihnNhQWPEd/GXn3iTRqfcRAVdIjuSjPvpmtwezS+0SBv+THgqUcAN
c/mT8VF7t922ME1c/9WSDuucVxGnP9PcVxxWwIB+2T8U4OyISXWAQIij4/qbJqFxOTZ64/lm8vhI
hJQgNCy/RKaIRq/dQ8/arB0oFIzf3wcIUyx4FGfOE9a1Vrz/1d0KTYcYd1dlcLEIrkvKMpuqHbO/
6xTW55tv2wxYvne8qiHGxiTk8YC6EW07Mk2/Ettlttlu6YejQQZXAOHh88KAnh0BzKpAr4Ik89kQ
KAhtVNyNbIqt8rVZZbsfBx6+5roiDbjI5anzmmulT99BMB1QQQAujvYLSvXDAE+dOgi26D1MnzQB
htKm0nX2TMk0BFsb8PHBhoJt5giKcYWYVEmJGsk1eY+vFf/H5avXRmRlys09NGf831+TUPl7fy5t
NIjGl8cAp2JL949w88Tondnwx9EMaticc/prOMfnzQHXbIq6gQDwHS1xUOeTxLZbTlt0lk8OVCH6
5TieRxoSaF73VtKasspMq/43kdXi7X+0NzKOjbaqAp5TtRR9ND0yULXPPXxWm8DCyXjbcRPAb6AD
J32VSJNxHKcJdw3hAXRO8KhMKzkDs+cKAd8zF+tFj+JHbf8M6HWKqoIrakgOFKgYkAYWQSNxS1QK
2YIQGV/gnNk30t1o9zWChCJQ7k5+CyyBtycgKQcAqigVHDKrN9sW5on+gfZ2iJeRqmkLEk7tKRFL
iOGBSVY3+RtYjOtaCyOhVOYOuhIXJb3b4QdnCfW3390bBZoQcU3mzRiUbJ73mFuInnSkEtKq8SFx
Xxa3GhYxBUxndqenFHFyc0o76K1U6bO8uXML5pWN7Pe/gh3yGIUeKksaGD6T/lDeJi9Vrh+ikAf3
vMXT6pVOMj5T9PVEOZvfHyM3QVs0ruCV1Q/XlE2FwY/bCh9VDOn90n8ilEM8uTEhQH4IwySgp2NX
hEagY9CJI8DmWDhBjKImtCIHg7g3kJU6wydlKGkx2ZjpbM6y7YjC012tDdDEPq45JEqUilSE8uS4
ATADo2So3OQpGsJwsL/Mg7Ie3gbEhRVB+bRXIDm0B25zKWgBRlT1hFGce5Ia0nsPa06MbOrD8tff
Ehlo/miR65oG8aPQnmHAld+X5Uhamu/6rysRazxkroVlQv9GiJ8+WRGVsp7d0wQZ0XlF+Pd7ucFX
OPIATrDy3q0RPmtmVAdi/itoyAnj7l4kdT5XxI507o2mIuDYk9uROiB8dBSWmQqs1nrfw1tEyDBW
ATMIHWY3wTkbh4sfQheO/boGj1TYGP26LrMPPdmNkSgqiFuo4eppI+Yii5rlWYR7oX6b4E3YGzX0
OxkkOQ2dqaz2QtoU8mZ52Ux6pHq4M1MBVWP89u2zIPF2Blm1wuSR+p6vrdXpCIHaY122uSSJrdbE
ajH3hNz00blq0QjBieW3YaZqr1EPVCnzB+15xSk5AQ/QoxTxASGn3S3UxPjD3BSh9SHpts3nUD7R
8nDUXn7sxfwydhQJnQ3BDh0ovZx4GnYTZf4Yk2Qd+ElN7Np55FilDI2ERoi4kQe19aIp1L1G8FLB
FmQmkOfauNjFGdsE0rRsphABfl3s0AvneYNf+uGB0rMhytl5lObFici4L/qvuQ61DHnuwk6+oea3
H8UO2VN6yLdFAW18+jgzp2P4WrjlFeIJti+4FoIgBxxshxv9EV4naxCnT5ak1QqdqYrVMOEzgvg+
7rpm1dvUQ2izXiG8/XSAClgPjfwo71p5eZhExFnp3x/mCe/FUSNhhKxL0VEwigZeJjPjrnokrhkO
pCzVofm4kkSRGs3UoiF/3AdEyPSn8vBSUktL9njC17jULr/q0kbescttt7lCR+NgFmVOdI65OKEx
XjROOhoOy0KodBIStbgnVE0bWDnQzQacpakkGgs73sGDZ012yMg5aySMSox8XQARntRpggtOmhYn
INV7d6nCxEyJDo1kkIbzjDpBhRxDkKpKvV/VUXr/G0sK4U/lwtE63zfkWS6Qes1nm+XeOQAehT1D
16wPYToc7c0nXhx6kEo+X7HJM7twb1YvnDYBnZQsBJ9/GVsnhOSX6A/POepd8tOOdXF8EZYV/TZX
ty4lv8vsBZ54WtiYIhV8gCSZoco3p3q+IkI/9OBE95bXnZHfEtqB7YDna7vgpnMRmHmDDTaTDW5V
boMBfLJ6p6TDNS2ULAG7QhNi3SK/oBSm5in/gBlcBL3NmO8r34jVY+8fcdayccX43AVrE/udotk3
irpdyqGdF5g85CcCONiyTrWDv6v3utT37Kxam3p+W9pyNSBfrnFo+cAafsaW6mquphtvzdp43Wf2
SQi72pRElPrxa+9kcEnA6JvQT3KLnQc8IvZCFHY7Xn7XHaI/erPW+0Si5YVDaBt6GjRkcAvwfuso
fndbEciDwPOeNUQJF+qLedbr0gYQlVu0brVUmO3JoJv5FPTUK1Z717YnY3wGyoCGJfB7LxIoivgk
yAXv0OS53eeuc4apkAHcBQtJGePtqcMDoM8APF5x30xxMXWX8iAtcCCddHbrinUm7HwVjFNBNZLM
/+a9tDIz2JfzE53LHIGy66geunGBpISoJtZQcmK0heOCL7gc07IvByWSSwoxf4e3rHwEL5mV4Ehf
eWJwc2GOL3ISp2y6+wa3HGPtUvZpPU4CemwL3c5nxK4TSycrTBP3Q74EGQ4iQlhb4Pqfz96Dbn1o
weNu3/MoAxhJ2LKTMqQxbmGvrcgHEwphR32dxjo+YMLQawN8qeZGJwBLwjrx7hmBe06NJf97gy0N
4a+Nyx7+sGmosN8zmN4eVNYLsU5BHx6HJJPIi/+OjHf6wBzgqfwzRLX2Qnd6QIvqi9zHOD5SQnU1
269C8wRklix6UmCx3+MxeCCUzzHyvaSc8olrk+gMGLrAIPrfcyiFrQrHQ2LJdSsJ56arSZpsG2Db
GdnzRBYsEvWPNG0pN1Mw0rrOC0VMmuZ3SMEEdkrFacb2gwxScymKp786KKnIIlBrzQvA9Ql1rg3d
AiS07oRfhxOOYYhWgRKCkv1HmDj7c8y0dfovRzPum+hXYNnBFMIz7aaLQLkScrRl7+EiW+u66eOV
j3htynnpedk+y12+7ABUmIqs3FaTnIic9F164TDWGZgVjy8pJx6YayHaoLSTd+yRLw80xGeLZScB
aBcKYIE+OLt4+yzwVmJrZw28WgV4hebVIsYhG9ggvfhGtFJSn8AHjcp7IKv2ZfzMWNaw3frBzNHM
S6WZ7dfqNZWzOFLCuT6Afvn2bpSYNic0HQ2CjwtW0V+yhYxocd1WQHCrSIpQjshB7u4sPAgRhUdI
ON2wLWh7eipCF99w0LLR905nNAJVnhUIXMtFko6dfjnm4iQnq2KC37c8et+hskMbWSQ43hKET6i1
pESYn+lzDOgVgxLdK8uZ/qb6QXxeb7spgrfbruFhTeYRhhP4PTn2fEfN9ECxZhhRmKBN8wf6hY6B
m5nwT9e830rw9nzNYXdu2gtCkXw8GsVFMKfqKwB0bktT5tLA9aEsh/bLHvIvhlhZpI85qzdE+PY3
xpWkBUFwdljKOGZU8Eokl4XAxWIbnktCd28peqoRLFU4k1KxtjRXVAKsQDY441lSiDU9I5ODLTTc
XQsXMZlXGra8T85EK/R82gsaURgbgwVb1bIHRzi7j3HEb8Rrkpg5JmX5J29B6qh0XrOhLqPDQXF/
1WPD4M7H6r+xV/qsBZMBW34nWwMUIJGZadGWEWwvE3i2etNprHrrBEumBi4SF27RMuxpHJAGAj8J
V79rYRjVQZo3BsmQvgZwITUQBkM5xilLNSzozxKZdNDXKQTr5Bt5Fp7DNWx1P7LiqZAzvvlB8klE
QjdhZABPnjG+QVkvLnKX/3lBhiJXenBsdT9AWfaKzvJgTA/T1bYjUhOuGAp979xKYb83QGPCamgp
HeSXlLH7f+Ib+iHhIJLiTjgRsxho4fDFmUVpXcHsg0ZEYY/yK0p50KoEszjtqNCYt59ZjMlUNeDt
uDRJXRe5rJ8DrmiQH2hKEd5miU+EMsQYN/GoN8mOXsxtbvvdG+ec4npjAWpcTQhX/h33MZv9PTtS
fgSXr7XxmcLnhPuP0ThjmhMaZe8ZEahYSSNnsWq8qR70SvN7G44h+KH5vgBYS1StMhfoJ9RXnz2h
IuwKR0OsOiod9T1KhQyiO+T7NdVbMIzEvqGUgOP9y4GmkA/04RFwmR/fkx4YkP5s7coAAK7FnhHP
gsPONenpsu1QsQwIwADM6KkiyI+iUfqP190BKtzceu9Zn0HZ+pqAT7VIjIzDd6kN/xSxV3pUjOje
rlKg9tRWQunac1ogmRbeBKiRrcy6IwUlcfv0jerZd0k6+gUDhTR585yaUev1O3jOMYotxQU/g6QN
cVvKiFrJoMx4T/YvH2nBq/pEmknv5gsY5ECMXDL26dcAM/TTJObPThrKFp8R4AJ99pydy2p60EM4
nDI2Zr4nCgPiB5vZ5YP8fGxj2XLqnYBzsnhqGqddyIBGQpKCDeme4crh4Eos7tyQpzOkDkK+WVos
aGzCEZM/Bx9z6CWe/0BOZBKTpKLjyJhZ9rrjkZR8uJvXiOpK7jVWj24F0wocwZgIQWnRSC6MJYVe
HXeqFvqCj/Ok/UNsJTPYQg/pZ8qysMAFnGy2FPEAvOaGS2Pqi9gZrfP/vIa4dkxrXjdj9YfWWaq5
qCFCww8itR4GByPpsw2YrkCbqidmDIZneAUu59Erls6gK3ZnGM7fX3/a1zFol/yJod2IZity102X
OBvMsp/s7DkmGJqh0RAh0BpejGEI6dUD84Zvg5fb+0jfTI5liqKWtMsWEcYHbxPk66SQbIqW2QMm
omedxNujADgKQLud4zj6RxBKdOIetkxw6txY/hCNBf1mlTTQHL1se6twL662SEmQR/KJb8w392Oi
m2eV0VXlbSsBVjSTPy++LKGBvg2SRTf1SbXF4qSgHskCQaH2e7KWv5rZl9ZRvCeOEq+n2pH2B1d1
kyhC3a9Em0LVrDU8ZXPNFvVzTSItVdlPwT2r4FW6nRcgT7L4gNV1nIzAMHVSyERxPxUsP5/HRSY7
lN5nVwEiA/+4RQL3aiZz0G0Q95xDX+SWTEoJpbFLXGWhcX7BlA5lubx8lHKMeJSBXcmKdM6k4NIy
A1sLGxgZp20qwc7cFT4M8ftT3XhV1wUzg06ooBoi0Ub06B21bGNLudERBsDwsGEvAOZsT8CguwBR
6iEK5r4phQrvnaPdnOKWssMTXB2Qsdu+7kAVGCK5eRm2GuxKQT2n2KgFKDT4vgDbhiZLZ+UDpxPZ
JfXD6+G9Wly6WBFTUjwf85Gpem/vBDFdIcwA8E3FBIkI2DxnhGXErFqJY7JZhtgxUdyX/2qlN76f
DUhLgVgEPWkse+skkjb5DwU9msHVegB4di96kpVIuuvOahQ72zYamABQvEalATalC1qNaEVNNy2v
cNOl4c1vj9PaN9z8sW6mwS3odIyX3eDoRbTMT9pQarc2gDAc+5DP7m2FAaWV9fANdvs78Cfjk5cY
1FMUj3Hzn1YDR+Bf25upESX335dFYouASme03+66u3CkNifMcEPYhf0K7rEN1jFKJWGA9H4iqZrw
at4NzOBG6LKoeUAQswQCQeGHDp930js+U7xnomm8mJLqCYqEaNTTgJ1h+yyR1PG1kpzgSTbzdnvO
JQiH0vJNtZQ6M2WBTzoOdLHtfC1fmkg7IqfJEjYsSDL8nkEcF6pHWO7ZbZDnQarCKka/f7FXpMyi
tgUMX/8DT9DpMqUSJri2jAAaJhnORjh07b/KrjO3KYIYEV0ttBkr24yCogFNKR8lmwpfs9SB70nH
pILVB3biyQlas6QwUJ2i0u6tGaCEui/KYvZ2nrW3HgUsn6gZH9GRBCAen0B3UEp59cwZZk3mrCk6
ZK91jdkW5I+sX7EKNv/gfX+rpf4RGqxQWmLnbXEGBcJtu6nUoO4XbIeybON0udEnyvMnR08cRYZ+
OIzQQTWhC2RiVNt9SRozMepmdLyiPTbQpswq5uczN5ElG7YidqyhdEuEWGjRzt36tLe1Bej44PDW
sVyh799iaLCVhbonQEnO9X5CbnrJzJ9S6j1U7X0dGbyZ2y/eBQDi/vsDlxnprkLC1B3V5CvVQhDJ
9jf1DLxr54ICD6+es+iB9xPBMUzmD/fQVyYns9gpUJPUjSG7AgwiEi2xeN03DO3By+c6MB/UyUjo
9+nSxkPSPQBKhZ5OosKczv+Y5j8D1iJYzh2KwqjBgeGP2Zf4WIiHyQUqzt464paf8gdS5M23iZ5M
ZB5XXXfl78a8Ae2TNdyjgoDw0mdS5cNYufKP4SUdqOjT0NZfwIeg1b+KS1xgXXzUS4ik4TgulBCu
O6+Inw5lUyiTC6fECr9Mvlk0yXKMzDPVzvz/TXcNDoiPVF7WgYAdB5mp/zL6fJOvTTY+r19IsRt6
UWnwDstd+NiW1ALl93hAZwsL4T9e3C90F6nh3GrhLb2f1f/UWzBDSZskef2QyYs9na7TtGrSS0An
H9QlWrIVsRVlS/UmBxkJb7si5ca8hK7NXYbSS3ZdSeBhYcjbShBmvBICj5iIOzfZBam3V+H4e87J
+qDTWyVw6f1YVpTmusCEmkzmLsQN2pPlBIoIBuU36yV2CAzFVDRfBZ7vkpxfxM2SofoaEx5ZGLov
TzXf6dghmABor+yWY4RVEEp1x+qG0sKZ43c3GJXHow0+D82CpY2DnVxnJWn+WJGZbp3nOSiHetmb
hv8GGLWgYhsN63NYvnfPXWbdvhSxigJlYQihRDe4iM3LA9tSXgvbeVhfsePjc9zNbxu7o6k6WFqL
YqYCBUoUJWNlBIl5oZFkHkhD8ikl9q6zRtdXSzFBbD+Nof4ATkiCXXa2DUyT3lbXuv8NM7+TXulk
La4WZxwwxgHENrs16rHzS2s5U5NSL24/95Z2/xKM2uBCbu1pEPCaOEe8xB8BYgVOTqhQEKbSUcdc
pyLNAdTeCU+uYWmHPeHTtEhLYp5d3DahDoBNnMXe0O6PytUkSn5nQfAJ6ve8mKgmYTCA3RNYasOD
ixzP7haCn26VJZu5d3ierPGx/+0oIC6U6OId4A7w3z/UjZVWtNsEGamyBpqvVNebOHQY3RM+SGVy
GTec7HqsHEZfG9qNxqZi7Gx5T+y+4YF8JLFIQtdmV9wUINk9ga2cPK9SuvU5dizPBFK7BDJMeMtF
B0LD7wG4/+LWu7ewkYmffdwdxge0x8OSV5F/s3JvxEH8JC86guwdxqgWVStU/q/Z13y8lP8oMHC5
zM5ey3DcbqFwCoCUcyagFIwcRJ+Ypm6jpjEFC5nUtXi6XXYcjTDIWLHBslZpyLw79waT6Ny+ydq9
mPJXBIr51NHKhFx3iz1IlGVh8MhRBjIY/E4ykCIUOmhge2S97PjqhPYm6x0F2Z3SlNueQQ1Np1vF
3dQJwmzw4CVyBYAKanRvDkq68KgVtAiVlLQ1rCZuMbsfOE+ppRdCO7ivzjRvFaB7kV5DkIc2L9ck
BxfYj5jw2/ZaLvsNub85CRVaQWjSm/CKKdnVKwuY1Rm/JGeLrFeQcy3rQTqo/vNDTovjIJBe7sx1
I+poS3XjPnOBS5G3Fus1gGzwqSiCpD04shHgrYrLckcDfLtvWS7g2GmcChbOUrhMmA+PTi4DXENi
qe9GvAu7e0qnl0bLN5Oy55CpkskB4E6+zuAt0heJ6OB0KpKxGqxLHzudDAAQmjyAriHn/PIPYMNC
XLc5VsurNnRVG517i0TzRrM7hUYphX86yTFdJDaA4+BCmNWAUWO6NC+fV5waxZyQz0sWh1OxmcT+
38XVdDrvt233TuPSAo7UrFcsOIs3qv/R2eSRhzdyPENoXYCrCIMXqzp3/mThzJq3wN/749sE401O
zmrdtyd4tx6CDoI4LFGDuMxO3ZC4tP3lkcciOuyC2SEtkfKvbIdDFeUoPTw8HGI0S+lFFX8ezSX6
phzYmsi+dp5Bdpov5YczKixxqJulyNI11zjFie2OAvA2/JgNeLBaWupRWHBVYzs2Z2dEiez7Td7X
wA/BT6vRIL3SkNpfESZOKVr/O59aox6WMWZr9LhErNmZKVUTSM20Wpxeo69ZS7l1cLyoydiA1z01
LxoFMqw2Mt32qiwRyttk5c7VEcoI7jz8loO2l1ZJL78+KafaQbOiyo/alF5msfFBUKuAD/jxJv2A
qpNr0tlBVNawOWgdyRFSCTdCdM4w6jMqzcDd/2AN69mIlx53qIFDui58H5UMWXvPa8C7YICvtEdw
phmwRnAypoDiBHhBIUgDWgbiKI5FA+RemFO29OFIbS6h/5pZrB8NnVix7zwcBMb0j743nAe5IBAD
ooHTotkb7ncmz7G5ctk38Qy+o6Qk2GORZ8zMKJYkJY93e09cDKgzECxoJLJ1ujHiWSAKidHXFhOv
ZJH5iiJbbmo31UQap4/afp2fHYaK8AkTrWETKVAH7S3OCY6Rm/jEKPj0aYJ23fAO3R1SxXco42z3
AlPOcs60uFlnlrvtpCCKDQbk1BavodFRFxnODStPzux1u8cC5IW2zD2Nl2Tnmz45MnEJBAfJC9kU
B9bfuxoooGSwKEZJz01xKfiX9V/3h1ecel66c14nIYRU2B4KOwU21IkQVyptdILGAaEBMMmrG50a
5ly8y6ELAhkS1p73Nfr7AdvdAQ8yBOOxcoEBiHooy+pJa+m1s4esi/VFFuYMnwzJVvPdwJij+heL
KMLJtyzVMGCtfzC1tocG31bjTAGaMl7G67xvqtBhpyBFZI3uHhKi0fKfm5cl3TbFa+G/5dxgZpPt
Cyji5yiMbk1QeBONtSkrpIDjgLto4schA/KRhur1jaVMoSPACRBn7KwOGb03p+wlgC7IHuam07eA
RjSqLbNyPYX+sbpgV94/N78m7zmXuFoxxkT7Uy5kHzie21CGOk87bkL/lkEIsoZhvpyBP6PitpVQ
5Fb5oG4zIoyojqpXgjzCtrlXLKPScBYTI0yIy/J6KoBAkzDbJ+GCRTQs29FenQUKL/o6GGi2U/pb
vUEN91o16pIDbmAeeGbZlsPuOmDrRKKcqcez+VUSKghh1SRi83NQvbRnNILS5hnNKwoeDAuWdVxu
EnysoesQdz0ng7Hl0M0ubAP3NKZf6QHc3ruNc3R/xhOAhjcEtsax9bxCqvCJb9hP/78+fKCUrnPf
YCa7tCf6D5950XT6nYUOxpbeGyAEW3j1lJ8aFJ82SdmVjmbYb5ZarkVoqKnzgMcXW5O66mXwCppB
i9ldArBMAO0TvPlNgvzmKslkWqM/s+y3GKUbZGcyiVSEyA7XX+LxH6z3CDpSKa8gf++9HQKJlyHg
4kFApV0qjchRJvQH+YYT2F8HzWFIL+RV2XUIEAzbNiFENF4f7q4MV9gAiopFVzRD9ObxYnFEJ1MP
bLhJiTkLEzhiL8xka98sBPooT0cgSNiehwyIRwJPhDBL5JgSQ3tqLcnYGxGqunnXA6d546yQmDYo
w+cypL3lSal6G1e6LyLHP92mtE3gz+zWvLRUzdg+o098cmg26TO1FmtDkCfy0JnUUWM1B/34BtUk
1t2YpGnmjOvo9NDfz+wgRqa7xxrzI8irJPdvg6Ww6izOhxNM7voqiGQHM75BbORvE6yCJ+m5/YNX
k44Z4g1O2MRccyCcky3KBocIxXmTuK4xg5bnSkgrxNzO18GN9GYu8CbTn/kQzD6uHipYkXEf3/qS
8P4dDWJtMsIsrqT+LmoCmoZgFVJ820fXso+qb8Eol7pGJaJPpu4xCKA/LeJyZJYWXUgbtmyJ/a8E
uUo3OMldSkR+GQf9s0aTSapnPXTN8tADH/R6T6LmulyGB88yzPsJlKK0bMMFgYplcxqdm3DWNZ0o
u5bQj7BSE5ncvXqdMe57H9+HZJ+58X1iOXsqaFfNY+esNAcwKZjKIjQWvipWQtEXEpyWlaoz7zOP
03QNQ+YWQjNvvb2nQNLw09+65+EMYxvQxNDKQjQ6oBohwOpa06ITPhxuXoV+b4TC/0IATG36ncTO
KBU0k2UiHNWdXaJPwdogglmCUXnc5K3vFaG0xIpn52j9f0xxMIOCvFWyk6tCr8FHh/jOqXLJX/MK
jx1KleOdWKD/88fKvdOwX87H6cBYT8mz3TOdh+JSM78w19kmW3TDy1NCwCYKhIpK1RPhcJcgxjH3
EzyKM3vtGELFRzl15+6A4Ji0tL1+9cAxtTx863n8mDsKywQlOQkwMpcsqPsm+ZlUP7mdp3Fs7Ojm
Exm/UtOoGCV3SmnGVhYY1En7qqxCsFTBmDTBOj+oNCe0qpiE5skTWLDN8v7d12L2rVaKGKgRhpbf
87p5tYqwjlPHDpa9zdNtECCvxsBlpZ3fvszz9p1KeZTZ/iVIrheK7/4dZInMeK4DyVMA5nH4u31K
ew1tITmxMluYIKekRdyrn7LW46sWucF4+R9fuTt5ZC8yMbEWAAcnkC5ry9p32JLGFiIPqUGQLHgs
d5/L4DzEDzbM5zSF9iSaVuzDaL9aW2CJcydE3pxrPg9DfJaH71V5tzElCQonQsJk96lKTrfj2sg7
98BrkjYoZ6RxM10s7OR0fyYRu/h+6+el8KPLSr1bcfx/QrG2xCw6Wdj3OoF06YWCNGFJdxNzNnrA
L/Z0984DJnRNU2kkQZT+zoUfGkdVUodO0M1GvLbMAYpN4YyrVCmMXCxPPTG4EgkyVndZPzPxSK00
fQqfqjdwyhb6NFekNGKZFDnCsIsmcZzHDm+N1u+GIdjby+ZIvokVN1XLhqpRsMItaTy7Qbhu/A+K
p3t8mhkz9dldPDzJfktuHnwsUoLK9an7/npxxm6Rhrb7peRdb4xlMSMDxNhR49VHgzkD3dAFWX2M
H1BxmMa6No5RER8T7DpLNYgGwf8u49AZEwv7Ia6vbEM2kN94RzebBxuXwqYy0QwUv0LeKZY3IvKu
z3ETrc9B/xJIglMLnSXSPuNUcN0B54H+8J1mZWyYKyYtk0mmeXSSGG7tdGU8SLANMLw1Ln4/VqSY
nerGzLL4AJmFPzOUVOYJWKk7KjehCw4d+HjTAf7S0rPptF8euQCGZvZ3Dys2jVXZZGte5BTeP2De
oQp8NV8rLGDN7eKVqHqthyW4fOI7AMurnPVxmIS2JwZB6MgRJIOm1nsPm6VJB6gJEl/ywSoBrPnp
UT57Gy6MmWWHAYS+YZy49WLgb9gdN3aeNCB9nX22eI8U1VcVrlcUPMsDt0v67ZwXBvIocmk09lFv
2cAX/OontGwRnFQVyDtYoNIbGt4Nyn22RbBGjN9TL0lQkhTU81VpHspmniCiIL52xWKVjq6NlgFm
rCthcO048MLmO1bBf/2Wqeb6T9TWZDe7Bt6SOo5t4/puEy5y9hmjicSFWJzs5keVIB5pWODz1yN0
2tkRxMuwsWuKW8qC1vXAKOv9eKG1GC7oNsjeX8tTcD1E2jFUo7eMTFVE8eiDTGjG7Y4DdTowd6sv
BpZES4rtykHppttz/ee6M7Hvrlp6GwAyctERLfkb/beWrUpQy96KuOOEbXoz/cdyzuCmoYW5htTw
C/CQmZ/koHP75cBp8TV4SKo0Tapi8++mvq6vwDzCzgOj1ShLG3u2BmwT6KBU6Ji98bS0LeftvP36
8xiSJZm2SGwobeWV6FAOsELZR61DyqPz1ZqEd1RqgWB9JR8a2NA1C2raRLwRrg1KS+xCCCLD60cd
z6+zTWwiG+IizIA/1niMdZw/kOx9NVQX9OdQusR7SVMrZGsr+IVx/iSMfBv3P+CvgfMzQTxrZgwI
F/f09sDYh2sD2mksj9ibI354ne6DRwvLjK8A59PI+O9uxCZxwOqyHqsYY2/U21X5rE0mg6y8NGr8
HmFZOtJcSnKtkGRpv7YoTrgxFJZoxiLaHyLiuTb0p3qhwiuxl58fCy+mfozvSqCEQ7BCqeH15vhL
Qk7fFs0C2ghzL9j3N1kJJ4almiKY1uatxpECKdnpMbqVwql41WbpSxndt7EiY9tHDYATcGYd1yl5
q/jdIteY4P2gS4X2puy/qN/IeW9NXeJhl59lnUn6ESVZ7yiURExBN8VRZSc6PjVITtNeJQFXVc+3
KYMkWwuuHj1691FGwk3QjtUkRU2eI7ep2dRwb1ehUf5YuB8el5IAt5BFBWSyu0dqui0zEppE0Lox
HqUX1+o60T25nPASwQknjauZ6G6rUXBtq+66Ni2WfgEl2ZLIDSp06z/sM2RvC1D1NwjO1IlIdoiE
HLIuvtVg3awZx/QVqSEcTve7LNVZP1IXtGMW23snVlp/1Oo+TkLYGmnmwEG7JGpP5bBchPl856U/
I4lUtYP/lvMKeBlmornvzKfxvPEo4hXP583N44xis2PWRuRWBI98yRcKBpoHs4+Yprqiv/ffjLUm
x+XwGpjp5wXYH0VYeyxY5XAwiOlJa1ofy1z86+V/xiAA3samyKRHAehWmAyDhpnQBJ67SRvQfR8D
b5bru6EWEC/FtJ1BBzb+ByTtOewwlJ21k7ch0ilQoisSInEhKpb6rDIibdTOpT/w3GEIpFjV8t0E
BAFZjACo8edwSMFMH5bbTzk82V6K66GneI7TbBv62Qk+8+9DFc2+WVRo0VoTjqGyeypRl+3/ByD4
G/jOypXIS1V6KKygfUm53Uwnhz4mYQ7/wIf8RScWSd7oHDOgzZyoboTfHFtBYQ5atxrb9sLfZ4v6
NvD77PpZ2I3YMPP5uZEK8N7AAQn9nVMTbsLOoR81LqMZ12H5gBHJFIIASSXdvjywfK7ZMcSzDncI
SAMTEpnX8KfE9qzERQPvhYtK1vj9dbPIdAVHmGXJcJ7iqxoIMhRbxarsTESNLayrCpTXR7v/OWhr
oeDnzwLKTlutjBRiCRTURCBt6v4IyUzXc2478oxhc3Z9pQLLqWQh3VVFzhyOwk7C1leSnuYfs+IS
P3ZM7Yex/AiZYx+1aqPWS+RsP59ED14v6X9oihBnVK3gtXtdzFNvr3y17IvzmGNmB3VDcs+AvYYZ
A34I7VMyQPt3tLut3KasPl+dSXk+Q/FMc22LxCWG/uBD163V7ipswAWtoBXk+uUqdB1sW8zWvNNk
p+o/oexhWyWlsC4DCfIV5jO11VD5sQ5wyzx0SLQIamtX/3cSJBxUUEEnWYrs200Ah6jdvYYHfDg9
bcHaQXIBhgxD6r0V90UBWNLQLoqLPrFMUkOhnkAicrZWS5ehlmznjq7X6HOmFbTl0Lmk8qng9beK
KVPX32FK/g1envJym4s+q2r0qOCmOhO1i0/g8rIYR+jiYVca121rZu8Z4QnW9ouYSJJZ0ooSg2u2
UdCbYBR3J5nMwPZMW2HeUwo1X4OZrEZHD4gdSzkSVS/8vVKuJvUFNyhMdHldmkOpJD7hAOof2uKA
qZ94Qs7RANyWVqLxfMo4jdvxiyZEEWIEtQyclyXFzNHv7+ACX+SxSGdtTCfaTj8uGwTLfgSdsi7v
cZibNoY15Ej3Rurg7oODELaoZfy5ETzmDaqbV3ghYNoOoI8z/TaYuvWnL5uzxxV4NOKe4QlcOQHl
E0g/j30XRf9Yj848igaCmipYM3nFcu6MVeyAgVFDWkfAi1dJzSDHnpDeZbX0qjBXKNNzMoVTP914
Tto3YG/wh49g8Qvxbnfj8Vm7uaJgUSuWyj3xbeEQqPMdaXSGtDMEp4Ap0IEOLGLRKK2sdtGa4LB2
zYLwHJSDfLuGykVaO0FX6tzJl7izOK0axBHFfs0C7UOqD91YNgWP7x9OFSKZL7x4eTAaxBCSTS8z
uypDZ69Dih88IXO70vbXQ5BkNKw9jyAaRFLuDUJ5JcVqYZRVx0NygSbOHxZVZ3odAU5ma1UqXtUI
qjM418QWAwZ55jX3W4Q1cj0z2W1CRfRFZmYOf2nvAjy263jl4orvW2NexszYlum2z/dcRHsDEjg0
oIWcZtotHx14+FAvchhW+ElmOeP311h+7kMmkjnJhpIrfBFiq8eriGJ/ho1Vsq8lpUcmf4jslqLS
qYT01wfagVNBI/OGha0SfCzv32MXTi3m7fCLY9mCaYdwAaO9Zh/fgTvE+/XDGAFxNxfUjoo9Ahjn
rHas5EuUV2RThRyR+C6VFRoH1DZTMTTh7x7LXnhUHYglouwnc6GfWYN52CdCGDsARvW6ZCqONKP1
45JBBAVs4DZWZ3rcuNE7/2HFAglMRcqegvK5nqM84H1nSaOHcKMoZYJpG5xibNSO5SEUv07puj5A
zn8xDEGOIOj/D0pW4dOWF4zhVmfeg8K95t4D+yRN2yZOgwdrZaAEKXw43VDcPKze6FkS7fSYUCVK
9Q3hwORDhpk8NveL7W91PqsnU42IRJvzZ43/sPpkGHNhER5MLUgTNcuqxAwJ5m02vCaVB52BIDqY
VydvLN9cNvItyboGAa8/5wgsHEPl9cjpnXZ359Cciqk+KOqZZkY49Kmi8tFcjpgNbHyrj/Vgaqr7
6W8YnachQsC0NHad1VcVn3J5EUd6hGQOHpmrcbnq2FW0qma0ai6LSdG+aAFLp6x/K5SSgZxXwp+9
fZgTV1cNpvlr1RiOJkiwqhIPwuY4tCF5tbm4BtdLxYDSNb2ixZxkt4DVWa1J2cYf3mQ1UV04yU1m
rw1KxLdiZ4+xXCDG4lJQYbW5LWdFo6H0ZH2av1oseP4V1a/p7CoXVbE42UvhsogPqyzmh+CmTmtw
/G0JJ1S/gQQxpnluGz6Wg4CKsVvywBs4rMraj8fuVoOdzbKBKS3puZPq+a3zjaoKZ3JI4VZW8T4P
iaXY/EySQxhJ5LOfpT75Kl2iflTMjinJStZj3BqDY6EBQOru4LByVU5XR6avDgYvGCL3I4+U70c7
s10Lmmu5sy3JmJZlBaD8oHwHEWWh0eRt5RVhNgOdoapPTN0XE+S99Wl7wYwB1yLg0Ik0ryeE1Qnq
W0ooFO8PfVeWVoj0Ex9JcLJ9IEvywmLRDLvf+DSMszpNLxeHukVis/QgtMqjt5BMPSPjplXosUne
XAm0YjTzhvK9UFSx7kUJIvmogI7jMI0tDmA1ZwddcTeFCI1i8+SXEnEYzfxw5b4W3Fwbyu4jWzg4
F7GV6wfvqcVqHiqNeLR1J4OALywdYmmwpcT8pup+LA+q/A53DkCeeUEdRnADVZE0c1ryHYWBSFRr
lKl15Z0VE/HUsZOnO48LmrjPQOxqOi8pqM+prFKVN/fl8oMyREOk8cQnmlIYKpHqxE3seuPmpPJ5
NW1h+J54GRsZa/r7B0dYA7Af8CTHPFa2/2BP9f0Y81BLi4ol+3oQskWlfevj1n3qHZdvIWoWCSLa
e9RnMOOrYbri8LKk8TlUoFR9/A2BA0an8hzgHhW/C7aOdlTuXq47iCwKvlb/jAkNoaFLDUy2CHMC
DsVOwKCclSmKZlkyVyGoWVoynuLrUI4EkXuGmncr2WD3jdJ94/cvycymx4lPX7/WDvE72taXhpER
9iv2sFmab9vGxGZJT06LCUN7VNEM27sd6rnLP4j9y4wmZpix5or+bYNCQBqh0DecSlaz+fiSmbDU
0dljVROptldUnEhzbRDtnQxDm0WpbFiJhzR8wn/1/J2xGEgq84DHzxX4Xz1NQruVcuKFkbXOVJg5
udMIQ8GAREREgyu7POzYRBuePPL/1LRQxiNI8sQZdsccSR8vCejI9KonWZZSIoDWQIGZozVmHf3J
w97qRoI+a+VOmkiL9w030R1mLyXSfa3fjc2LOIiJ9/HJhHzRTGoBpB6kftjEFkr522ys5Bj5LQgl
Nc7rD7c4MFGpsE2N+b6EoyrJNMbz46VhdkBtQ6lebuC9e8TknOIJAnWUkiMqTDC1pWMxgHmTEQvb
CjlhnaSAjpqenepecknsei/d/1TEl+pcPy8r/MnSE4ROhXW6IF+dMNYUallF1cGsNgEBxB0aZoku
1MhI58jHO2FD+gXGl6iECwAJTTcLTf+6X6j2NbMBBy9C32JJSnkI857eNgLCu+eV0y7n8FZqO2Di
Y8A20xU8pmWpceyRrXDOdYP1WY2tvvl4OXRyrc80omVwTbq0iRxTEPX8eje99hdKV9C2u8ddCWo8
EXkxKjb0xx+xzz71E2/5dnrPh6SPXHgV5pfyYXS7AesH2T9aC8F6LaalIKECDmq94dh5Ejksbh62
Nj1xaju1KyNP1qHTMTsnIF1Ahquq37UlyJA9TYf63bIgSZ1hooH2W3ksOxdu5+7/ZMWLH71DP3nn
c0RRd9aXdrIrimIgh99ldtq2eGOe2AxChrYn1Eylmc0cjvcHRtVXR8NX3m5yHBuDfphOxiB4POwd
Ee/bWDVUBmNA2o5JF7qRJ4A1+1GhYvzz4fxSzVRkP1UsvXw0XZHRKP6AUY4amsd0VaE6qUif7iNO
TRJk3Rsau6m4iBbuCd83ozVzCu/KvnRRLgZk/nUvim5a3PTN2KTS0gGWCVTm4HAc7G99q3ELDJ9R
2aoewWrexkTHpx6+fxdSfFbgPsGWt7Hm2G3rpcu9Eq6F0sthTCfmuQ96g3zApzh+bq9OkNZqV1yu
S0/m0hBbb3HaYcJkoZkB+4BiVm4v4M4HjE79P5sfsAwrDw0BLLP9xK38xJYiMXNmEsVGycNOgEOQ
E4s/9CbCd5Yz9Se14sWCoK30rKGehdGWWXOUFXk/NR9s3CKkrpWxwbgy2KhQtaC6zTPcKspRcWIv
NgKrELpLz8NsCdh5Y+aP9MxYSvXiShDuHxYngC9Nrtot6VZPIyFDpfaWmFRyoV/Oi0AM9oy6kQMG
8cKZzeBFMZkeoICgJpgSWNnPbvKrS/0YHmsT2nnszemwV+kK81t+zK9H0LlrMXFIW6AYSbI3dLwi
vK3s+ZWzpGnIHX4KIsPsnnEiSDPhq9Lml2yKss4QTxiw/2hRNs6Ex/3sPNb+65sjav5S5+begVcR
SzuDsDu3axZFgz7ZQyzMADGMgO/OVkzo9hP3V9p3J5NQuYuMZ/FBvmz4Mfzb0abdsN0p9JTk3kPA
P/vuvT1eZtCzWgZ5rqAGxPXokGxjVG8KOG+Jvffe9Qz0crt2Qb7I6aGEq6Ft0uBAqzAdZ+BG6gU6
cU41MybaZfHEZoaDIpS0Jxy650nQd+xDO+o0G5MFEN02DXQiuyRoSz1qKMsO5kmtUviwcmmbN9Ck
BwlYppZhPQmtnvdr2BcuEr7yr/6ZsBwhCL7iQLG3A2i6lJHlKdirTPI3f9SYq6ztHu7N9xdxeh7W
3BXZdzCcPg4dfivEK/ZfM5xld7j7tTwrpEIw/f+Xf02AqmiKYwoGz1hgFq71X43axFdaA4QGSAjk
KrxpcMmrkW/FyJMxgA4x/BR7EEpjt3VRzjEeyfwVtrnKpchLutrZ87ODzHRD7tzb9ZDIU9FHHRdf
YhsxH2DLT64nnYjCx33Jizc1i1HcyDqkt11DprxILPzb6ka/TkoZSckx1VDmO3IxLLepTAaROPL2
jISQtdNWpQfHIkpTcIKWnWtmRYeLS5XiuovKwYNKRTte5wFDyY7GZfaWZ2ljKyOYbO2n3xeKhHuk
pY0fjGpUBGQ/ym04ZQ9s6znLnepKuN80XhlzDEZ9AuyGhNBgTIvDPbGU21sxC6JD83qlXEOlv09h
X3FWcJME8gcygc+WJjWjzZRJpXHVuSxxngwXxc2L71Bb85MwCfz97t/c4USxMgJu1z+XG9Tv6M/u
g1iI7QESaZAEFS1wQYvfoXbQV6p7yT0p99Iua98yoTk+qdwTJ+hdhb+eSoLQpsQu+I0Eupugr7XS
OOxKnfwU7P5lep1HT1841WPj1+eE2lRGGOWlNvBgzXEM+YsWRXy9AnZ4+2xJSvJC/ySNs9j2flIw
oUBPgfBgnKnoWbfzk53twFfFzboBxuURt/HzJX3mIXAb6teFaP95i29tgaMZ0HFxJcMjUCAUQ5Tb
F1ptuRPFJazcpDWsUPnDkHhCw7bYNy4fViX4nSMohXnfNu2Fx3yTWq4L8LOg7NGmFuvYYSVlU9eK
j6gvHbm2tm4o/RZfYVKxyhozn0CEck6CoAwsiuUoPxC3cxIqZSobnIWOFuMlCWLQkF5W4E6sOog9
8SjHcu9YhYzd8zbU6vXI+jAKf+PaQPnhOf9GUx6GMonZkwRB74veN4ywnQEnTfYDMG87Xg7xzuJQ
7ky5+Rq8tAMc/AvnDp10eCtK4fRcdgdhU7OjKNT2pCzxozrSg/jDCEC8rltZQPw9T2PW50P1wN5J
E2v3c13Ifzffn2uWjsjLnh7P2GnlMM5oBW2kuzNbnxM4Mrcmk42+o2G/tSj0fNhcPKvMMfvw0BDd
HXdqgqXQM2hr6minfgjsoB3nyuSk+E8yOvOwulHtJ0i9iCjkiMPeJEIemwYl5YPqK9vnwNEwHnkA
H0pdSDDkglHUjaTdnOt2RD1ySstMl774CbMlxkXoOai3ZujoY8nOppd4uQTHQPZyeDwsPeHtREB/
Ixvsk1csCxAXO4nt/KTnBTN44qWn5zt9/1dRKFncklwx0k3kkVJAApCgTcfuwy4PKRNxaCn/f40e
omuI3v4IskY6ZS6yuouLxR60nDQfLBwNqOSZHjAx9AsjP7DGJR1U7y9lqWIiZI/A+8RBjbLB3P5d
3Gbthl0azwW0EWp+M7oNSeN2JRWabvfIs6nGCBr+EAC6tzQaLuY28t68OvpTc1jxm8Z5pbY+SJW4
DP04sGfK4UkLkFYX8y+c1kfQk8xSyY00jhKQjcgMtGZ6yn0hseDkBSOp5lK2SdgIodG2eAJdQbgB
9d0DLEHXn5HnFb3ma/0/H1KEDSxwmaFAGktqhQEFk3fc/LLWed0hdQ5xHXPN6iIDFO91WKIu5jWT
rZR4cQkZb/+okVmQmkHTf7/vBEbuN7KO8MmzIrLCwPHU+6VJz6HJWRwRaYhCj4arisBOIj+FQ0VD
qvxvBD7B5hurDS0Wcds2bAHB9snQoXw6hPspZRqa/L9vBepQUC9HZAacfLDo4NHlwbMr7sD4/x2O
m7/fgWd9OOR3JogQREYb1c69yYDc7nOJkOOBUuFRomdUzwmBLL02m61o5CDu2KY3GPtssep47ngV
WDYfmlJ3+XPJjU1l4vAKiOG7soQN+EToZHQ1hqsZAI9phSo1XbkRgvZDfa1EaWHpSL10+/a2/tIo
Wn4Fa0b9BRBhwWvwQox9yr7RL5LQSX1GR/oSP8dg1N/iL6tNvdo8olQTJlEQs2aeDr7HLYshxBH4
XnZ6M75R7IXvxpwFFD78ed1NbhEt3eyLYQXKK6zxZHU4Y/e+gwB5IwkjTlQTvtamwo7GqM3EYxTo
Y0UbWwowj6St13rHQdy/WEoJL1NwlLPeeEfVKPDcFCJPMT+JnYUzR/HFUKHh2WvMPO9qu5L4Cx0e
IXMC6kz6UXF38KkaM6GEPMpdQqBoaG6m6g32Cvz6qoGV5xaw+kaIukWfVRcw6blj2XDEeiO9gaUe
gkwP2Wt3ZKPIjMj71wRg79I7s1X2w7NgPmurhaSRVpObGyxw7hkboJ9g4ofAY6qkvFGrEmKIWCPD
pb5JizAYx26Fe/xs8iTrI2Uo0lkQSF30todX0TAS/DVRdk69z8ljS09f5HK8hTIBB5L7nVNIXdRd
liruAhNqo2DB5imYC9rICcA4C0CusNz38sNSJuHgK3GLSD61FPs9RTFbKusmiGeq4xUdRAHLR8tK
i2+AS1JiWpR7tMhLWVcZiraGAY5LX7SU1QVH3HdBqTxsI+PZ6JMAbdSMfh+glhLoBx5BCkWYcw/H
bz0ZcNbQcjbgtW8TO5y+nR7N3T4ahc52z91sAP29LXGQxZkr9lxokJ2rxdYOKgSJhK/LJUXPqpGc
k/T5jNCj4ES0Ato8pAqPJviDUlBRESJjZUGo2HXPUI00FwUf8lhzANCV2LSgFNeZOBwTk6B5T/Hm
izR431cqkZ9ROiT9qrX1fWLuv50sbYYC80l5nDgnlaNtoIhwQJiUaA1VPGDL95J30mBDu5cM3Z73
IsJ1W0sBh/A+CWmJs/KserLEGOU0T8pE/EroM1ilMWNbqgaP7gP8q/gr/gVcZtjnA2EVB3OxCiiJ
xA1g8RQJOHhQEHmXgfPMRiZH6gjj7OzmlLXFx/dzXUGKR98KmP+c9gf2Q8bsCkaKNyzkzutIDZ9s
VHeHZo0Sx6JsavVu/2cZDF4mr5+8YGJwVgugqxzUi4y6wLrVZU+sn5y9qFCiylFk0RUbiMKCcC/t
KJ77RZvK1+ON8qkVTsCU/DVl3bcCzos7G/g/XNH7ogMtXAkUEGMl+sOo/XCvsWQmZphQBVqwUnKt
pjWmuD75LZ7S2Ha7WobcaoJSDDMzU3kPyXk6kY1cOCGjcpuEuNr87nX01bl/ZUXW76WEz6dZryn/
ttKwF0OGSJxyj5BvA5erOCO0iI5h31BIsn7Vz79q/bVdM9jyM1UU05lwdKI0bzFRNNo0s/V1nUXb
PTy9PIJfpo0rLYWZOZh0hFpJeMg/7lCu4JQoIqH1NnMWJrgsQGvCbFpkU8OIxJOh+c1hOqNZC91p
QwAPBHbWpJkuhBJXL2cArPkfUz8/UNcBds7ompKOz8mOQNFhd+R5tc40id2e10ARNWHhcmsYQAVo
FH8130NkjARp3XBnQ6H5cnhEw6Nhlx3WFnmssIjyns2I/skf6tjjPZhAGh1WRkD4c68RtVMQ9XCo
sXorZ5Mh1cmoSeZn7CyIT/K8Iva086/Zw3bYSX9tBuK4yzB9E8ALJM6bFp/mhNruVdrVCyKHMNBD
j//5tkwQT8Je5BtEE5bbKJIMvLOmSh9yZeX8hlihGkDMktP3cOVFKPYB2KYeMvK46riwH57m2VjB
PHwRIj54GYIT2LgTaB0PF9apSQ9Ah4AChoLUh6/Z9B3DpG8NLAMa86UhnLBJ00X7WOckmrsVsinU
hArBMn5/b3mAyJp/ZO2nFS/JLVoAXos2euuHR4aZ4qeFe6fFfhErh/5ipmXAGicvVLYICzJL2MBu
YFjfTBL91mdvoncfiBzdCUgR4wC0qneT4HmH9qT0T9cZdSGOmnuDKNB7AJyEbuP7vXclQSPbjW7T
Hc4R3I19pvrQeR3GqQv5K8zAMuZrcqU8BkESPtvHxw8Hk3u/35OF6mF7ijjdTtTNtoDEt5B3ihZH
yYvIWJK06t9VA62gmfsQI0n7pQK+FOWQFv99oKlcZ/dTCtlPQBG9Xox6tNdKb0hcm1ct3pomxnuJ
foyDnil83nvawYY7r0wSMCeohAaxK1QKpVrFnCVW+uqPtRgiFROWCoohlEuyCQxifCLM3v2PCo4i
yuyYA9dUPPqUHymXe2bISpfMN9b77hritHW6DOjz7oD4zl7yGXT5WrjKj9GcE2Ikil8iHkAUsYuz
VhfBrWED00diRIfnBCUxCrZYbpdZfRAUB42uuOhNBVylB57dVTCFk9+ZtlzfjxHhWHVRN7DfgzdH
pdECX0oNzv7KgTj5VGVtHfySK4E/oy8h/rD+tRa/rbLYJ+r2bqxyuedTUk8MdrJdBu8Z9j5LheDl
nN/YN1nNV4Ykc2ru+nPMa6/cb2/SY2LIhi8cg/f4UWJi+wIJPBgy/hqA0igUyIRsDH3pW85ZUDqy
tlLibO3hZKqyW1CGHTK4Eu3cvHjMoMQpH2vN8jM3OBt1kif4Oqf7WvTGZMyO6r/puiUUgn9DG1G3
i5TeiSCxdQUm8Pst6vs73JQ9oxLWpzPJeeLl5hqWUSmEgJ6fGf83ORDkk+g+0f0e21IakBj7eyX1
xDYjpryRRD4VNGMsqxEiKA5P6AoCWQExFrXdO3wtb59ieRvEbPRYUdrn7PX7xwKd3OsJuh+vYEyz
uXVdEdxGUKUx2iFzhR7onqkgaBRG9BPRJmt5pzedB1CciYNjI71zuY5xThotrLyPc2E7jdxhMZAV
+WJ6GG+yliF9Mp1PfrHdquezJskUFl1M04kxEKxu1eTr9fyYksRdhwCXZ/EzGyYmYLxmxG4Yl/vz
EKiyfQhKwxIjBnAgPkAZsWqHxkNWxj9eSv9uvOfPIUo/nKcQP4vmo6zWZcFInl8fP9qFsjT/k8fn
+cxVbUpNEcRCwpB1MO3QayE1rkAUeBSjZDuczhhZAdSR0hqyxGOrhfuGeDc/kfWcNilffrscGeU8
s3fHPHqKwXivOMnvHPVf2gSekm7B0vu3U+ROy+r+TKeY/LOX2/M9L2BMt+uNfcG+m+Erp69L8dKa
enja7OFUJTzbE49F8jbdfEIFhqBu9lnC9+FN/UkvKsR1gQ1Rrit8YOMivInZ2A4pZRDoCrd/fCtg
4OIX8uVIJGONlpkKBawiPYQfrXng8pt4y8Po6GnekP67XAA6ffo5KrXf1UDXl1krMdSeSyBvdDto
uXDGdnjtbHDbze9BU4I2u/oI16Ky7YPWBV5ODkUoq3duBV3hFff8C1/4WFULTB9bcTmEzR2OCcek
WIiX8f3dZj/xScmPHy+/zv8fWZMiut3tpgP8TouIOpq2MtBEQjoCOQi/rqzOIUISItYx9Jz3r0Ll
4JAm2PzOXvboG8kuP/+xstxYurs/5Vuy917HpQ44ftcRvvpKV7UjE/kyZlr++V1hiJBwedp0v1UF
t4Sx3xPmni6jCU68SIUuMoKcW4bQRor+Wh+VowWLDChvnjPihAZZI3+YTGbinBov72Wjb0irhdwU
6YSVU7aLnbHcooFf06snjsWubYRDXXW7BAIWv8mADJxvjx80cJAeIb/RhvASK3KYpAp+i/oXUOQl
jMAn3R9SH+HHpm0hBylkj1ml0Asw/T2qnO6HlFHCeykbAcHRif1OWrc8uSEhfOoZ7aXPum6+eOVY
ru1abYK7mzO77p9nMWp97MDx92DbtleZdixWMAXspol2iSKWTOG8ZvKlkeKoyfcGXlsLRG6evzPM
wVdi2050KVWuZ7HX3U0K3rWJmPnsjy2Dl9yll5GCpfCYW+usKQzEEBNjyBMU+l+J4c8MNXQwYH/S
EGrk50NWBdkiqzFFAqqycb7I59pvE8/tet6if51Btw9BIGwCS2TzPuonZEGxaQxkJXcFsjiybNIX
n4Ct9jANFBnbDfMFCBuasQ78osFjw5JK7r6gTgAS/52sccIwRDzyYOoQuUN4FooRRbSgO/Nq5SYr
eVBzPnTrPudsTe8FqHWL3yU4e3RjOvSyKjN5v9m9Y4o/e9EdR8OTnec0py1Wh9soxS+crcfCTaHe
HuQg6SISxRncguPrFFcLwibgflIcGUxz/dLPIPujFd6aKqk2IB5Nu+rECThakJarFG5stIgyup2Y
FYdz2Ku7LdgnfBHwMWDR6sJPrRkFSvSsHQf2lXo3PGRi+lAysfWZdTdPpow8ZJ983vGD7ocYTVDi
GueGKzyZGhwKpRn1VsV+uFFMzIk22VXXFCLW5mjeSJSfTQ1A5fDFDoyAheR7BYO/MeiX5DFRAMd8
vo666H8cQfxkPBbw3Ord5EUPKRMlIXSUUGo2cHNPTakwka8yjd0DlkDoFtiKJmGxfomGrp6Bi/p9
1QMH5ifz201x5z6gS7YzF0cLQL3E3vTHIm6EylmleOq8NAtGmHEFOnyqSVwphBZ4QZnfHTpvWQhD
3jvvzW33QRkMBnBqbU7UDao1mkgYC9vbnsl2DHTUuf53e3qHB3lHepz/U9SnqGEZYMfujag404p/
ZHYlJiRxWakbBol2KPl2rbow0UCeNyPdLaEVML2TOWgVJkd3lx3Wpd6dOiZN1cfKon7DgxpNJOtc
DCAY0m/70PXI/OqRjei3Mh2DABK/fDXZSIMSsU7PzUaRI4KM2US8ByUOICg5YZmTRpvtNSzFcYIe
uY9osXmtuCUXfeXsospzkDuIdWD070Hvfe9AD3YcBWA52G9Y4nM650ICTAohJ9+ZKHFFID5TBbq5
IhYWah3JnEI+gbjwc9AdQdyoq0ahlzhWiJ31CxkEeTylaRK35M7MfWPwVoYb7H8weKCc0TUARUun
TpzsWMXU5yUBhWBcqAnZUXy6oeFu0IzgwArpb7TULaist8tGoP+5XH14XNvsYTIp93jCDDOPVysj
Hz1kZCdwutU62in1Wj0W+EozCCns+aszUqYYtZSnkQtvaWxcSjFNmWOS9FW8OZWsrdCP6yLddjqo
sSh9TKHD4UnyTixkQoXsyyMa1Ycw9igTfIyV7nZHKpiNSdsslEmi8s9tNJi6Jhf6ZRnO05nG9tg9
e6xWIxqw0Nk+Dok0oPRH+5I8xzFJoa4ZhNTZRVipKYq+Y3pKVS9DFrEcfS+IOGbWVJdS3UnbHz5p
VU1Wt0uHON5ylJYVSxqp7/runHQmM33pFgAFKIbDuzhKSLDqATI/Oe0OSWXsn2Xq6oMHeKUX9fCG
eOLnCgLPTcZigUwtkD3nzgbwUA8o8uDEAHX3ga8OMcKBHOPxJSQdU3T+hzyPYIfbnmLAZ2t1vg7F
T+en3dTwRu+6pjBMcQ+xp8TqjHSCMzXWnlCT0zyae9QqeFuiNxU+Q3ScNKmM6k0iVr0i/GbAOS42
qkBp5UGZ8l6NY1Km7JNWaib2EV4xKiJi8hMdQpvCa2RZn8F+SOhuJf8ou++Y6q2MoayMGN/h/R4W
pyA5hOOyh+lKNczqb4rxUwKMCts9sN4GHGvEa6HtB/l4eU9/tziJWnJw99gCF5BRxKfONmA724Gs
Mj/wM7oJ/KKtl8LDMDusNLK2U2esnQUziALFXKI9hCU5G/2zsbRwR6q8QXAJrBqpW8fcrYQQBKKX
7mpao5y2tEn8Rg+jfO5SvO70h4gnJ8rvtH3uz7dDW5cwCj0kQP+eoALL2275J0HE9v8fgzZ0PiJr
Ak0dhTZ+L9OqYsYLjNqW8J512p7hnShSbP3jl7hdShdtMnbBhasFrhhfewceWv6k+eFq0JIjvzub
ZyYc9IJrHqrmKwatQMYZ1rz4vq5bjxaDq/TYooBYUO0qkAhYmh5TxThh91eDyYyLhW05rhVFhVpx
vQsKcM+T4yXSadiMLDqDY4xtU12FGoHpZllKC3VMnMGRKNowk/xWxRx5mbniMpGrdZnY9CqaPbRt
dSgqAonByaG+UISZxvvTngBSR+abgukWDximlBTG9ZDJe88fLTQKWlIpkruKsQYlG6FaCofWp1gu
KMid/b0IypBj4t2D0m77iMGC+UUF0mhco0xdXrdiaT8P02utWjzdILvo8Vk8X+wz7O8wuGS598vu
E7xAFbLGcQjcSXErT3/ZK4MYohkpYFcsx7MTmsNjHkcRvRJi2NfGXtC9XNIdLYVxiT2x47MgCOV3
bL5EvJXcwaB4EluwFVBqF0FzOjVppG0S573sHsBfI3lTit16QMYZxChJLthjXKCEQkpAVNjwm/Jd
E+kgpKMzCZ4zcaM4bsp8rCL3VenljRP0WEO7Wpv96MJx1a7icDZ1Nu6uc4I0A8tYmtRDuKjrQZPg
58DOg9k=
`protect end_protected
