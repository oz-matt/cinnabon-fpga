-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
K6SXbCNsfxMTrahmXVSL3eEjckVKmZ8g+WYa8WYqv0r//qiXnIjvGPsYE3b8Vr5wabQJtzdVMqeE
+2zRt4WVo1y3NpQaBeKWLSsskZp9+F0cFnqztOIycb4m1H20ROAD/QLLw9wCnco7LZmThCn7hdy7
fNjQJeC+dDA558dO814AQCZjPTPTYMp1j92O7jJRqB+VOHWM1UoZ75S4cuh1e2MOSrCaC9n95UFK
0fBnJO3l1WuVjMcl3EAvlHaYbnTos2OYB0Wqsh1pmKLT9Ug+rPe2irlFTbg1K1N976jjEfeeoK6C
6ilCCF6Lrh1ow7FVF+YOmijzzWkHghK1rhoCow==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28736)
`protect data_block
EbD2cUHiNIiOFiTHbFbfShuH8Ar0KpoTTwrxT7vnOZCJ6o6XGweqjc2nUsHQeyZ5+zdehqHwqLWZ
w3m7ObQruNsTThbI+V8Qt3BR1KCwwjO44lRV4vTo+ZmAXD3VPpuLOze6BIWygvxZ/moMuJOSeQhh
Ti1BiIeHn9NKOo4mwznqcoMm+AY955wkc3ShTnDK6rYJuh9e/JjDXlcI0U5A2WegELn4p/iHYMTs
pXNHt9PblfPB+cNRXPL9xAUy8aHY5cmXV8YR0pPiPQvdiAKjENui4+bbcbG7o4fRpqWTcYgXfb70
vYTzgnz2d6Gbdf62paBtT0c7Yekdo1p6kQZqNkbMFE88gqayAG4g4MYIk96llFFhF8Xug4UPrjsy
UiJuOFsxXmIuwFoQkGFrwW8iwM+5nAR6mxKPVBP6NcHrFB2b6PABd+BW4FUlogz8+oXqxRBoUHee
46IQWskvdwW3QO2khWfI0OEUv9fUZ9TJ3UfGrbB/tAnRR5+oGGWLfcd3qizHWfLI0Y7qn/o+94L5
oyYvxruWIhurGY5Zr+/ilpLviaKti1isRRXVBDJ2VCbbRLfI/gi9c3gaQ2/Gsru7Fq4VJGQKdD0H
butPK89/mbRxajpvggoaNf/ZlGqQoAVUpVD3veAvWNVLH+OtnsJr8Q92G+pVhGDyNb8O/fLTRsot
omhI/s3nGVWmOKB3AowYAzgy0jXFjsZsEQOJ95/vZUXdDdIqtLCrpgsIQ+gu/bikl3+RXlUhkyRC
cTkhofb6yktHmgWzCQe1VWnpp39rx2Xadi8Zvlx520bTXlLOLBu/ILTMqq+MKLxIL2KdkcYCUtpa
iDyso4kDqVN+qZ4dqE3GzWM9VDpvBv4DobVfVxrBJ2IdjH6FCksQFFCBhYZz214VYtm9oRDfCq0v
ULZO7n05qu4xb3xKfU7aUvvQHvddbx7jggtX7H6EvF8KThqubkTYvibVtH8DOpTfsmwKzJrJaiM2
RdQkMvhst8y5u1jmJCSKROi/yAZ2C9oL6VCNTGw0d4FoD+WH7mI/e6jWPdvACzP9jl4S/0EksNP1
zHrhHddglQOzrYgs3dwER31LRkN68tddWdQ9hnz4pQekHWTfqsiV3ZFSakM9Jc8x3O6S38l3ZuW9
+fY9faoadduuZkaejqvZNGGx7FzT2sMQOiC32tzXNNsrU3Ny+18N+HHOJBTLddOlONFJ8tmNSP4E
Mywmr4TLSZM9dwTUeMQ8xyGILRdd1jfvo8kUNu1tttFr8TeGLHP1ytIMSfdriKMEaMPLD7pEWqZa
wAxNwfwXZOYeLlckANEvmgXS2bz82UmjJaHprmJjEDPFT19P4Pbr1pfOAQNn57XSWsMKkbD8VBaS
2oJ6suThaxfTQxtZYED4u2p3iGbpKkflJ23hBaLbdQTea+QOTfT0W/1dVred6mezozG18ZkqyJ2e
JndGWwL5JbTqEnrY7aNpSmC9U3pudRJEMcTzTaeDg1bYTZFCx0uhu7AadkAPeg3FEadZE4xnWtdx
lJXIKtwMNKqfKrMjKJs+6tA/1DyMEA9W0zbCA40yzi+PDHwLqrPFRiO5VoW4JZCU0PwKwgK9p22/
bSTHxkZEDvk85u/1+utFlLfem80k154yyBIL3ER0O5q31ug6kHgPu+y3EviWYs9nqH+r9UGElV60
xk8jlwgfUDhUXLz3UJqfretvCaGwaMUJm6RNzWxFFJafTImNF7CVNH2nVSK76v+U9uUOh4tSkJ2i
/AAwk5MwXuHwBRsll00wlo2I2Sp4FNHjWZBVT3XQqGbEcNONdfCsEa3TtFWrzIQkBCPGg5lnuet4
1suSoC7non/vLMMSAVAK2Drr+svMCD4/yefwmGQrxzZBAJJU8M6lMOUln375Yz2A4O/0RQWVmSOf
PJAVg8P8m7CD/+0AWsgxxeVkgu/+lUcOYz/UfhEjQYD+XsRle5qmEIkXd4ZQP7Cm4ZO0artGiQkz
Un/t5v2LadQS8vxTGeUjzaMVNTEuTzcteY61Bt8GbJiniWtxBdS6g1VRTi0J5JrBgORtoBSbZ0En
GU4N1PBszsdCnxi03pYIhb4lOj2S07guToQmUgnqgIDabwPkjM0LjN9FAOHVr7tpk9KJa3OeG0Wg
NX6FfiShDLn0bY+3qn714MHrz0er0xTUi8/wcPYt0rCuVfVWv90jBLU9HCM1c36vkniRlRYxZ5ww
7ts6XzHIQ+/mPN4xhpKmIq6QkFJiXNPdLPPboRCdKSN8DhUTN7D3J1NAtrnxNq0hIqt1C94FkpEO
hDpHMC15tB1oIVJV0VuHLlzp7rH/4TraoIuoMeqqvaZOlLRr50nhBW4mfVligNU4FdM2vGkPIl9p
Vyr8fxTp3Z4dCywe6NTH57mZLVOm/Ppa6M1wbhUc0ZJCUSFG/OWTj6Dd/JefvkjbMnlTFnKDAiBQ
h772wlQhebtqWkbRrktU9aMMmpAm8SMBq46etdIDlU87Aj79qNJuBqenM9opzTqIAEgAj57QZ6XP
2AA+NEuD2HoRA0dHB/5ioBnAE+ZLxT8RUAzPJxvHbITnXd0TmiWcGJtxa+u+SbEgPox+8ZhYkf3D
fShADhAwo7xJKz5d2/b7l4DrbwkcxndvU/dZOyisG4z65BOSAAgT17J+5nHAvWTldnFnB8/0LHaL
tobrMzARZxbrrS241L7GOINIDYg8cvKdXuDAQT/HXGq3Bpr1XPJccUryMW2/TzMsxU0aTsjTGmtH
KvhGnJ8cMCR2HEdUhtiG+vEyvdnhw3cxlnoi9n4cQ8SPPo//oz1IKMhlokrbpheDrgVPWzvZo5Va
eVnv4sH8m+VzLA1rweqraYq2pXQfoW2b3vKMedJSezQp+2nlmCD6sQPZNL/t7W0699SNbMPXJiQr
7tiJ+zjibFd6BrSsqOAc824VqscbZvHUdR1Kyu0mHUAVakBBgbBt1KVcgE0l/z7A2+3h88Kmq/6z
HrIiSLVTJXaDsyRjYRANy82GB7+VZI59Q9XJzTP20NkO1QoskK2Rio4zIXjfdclNq0HTfZnNDE+c
QTUgr3qKGjqafPUqzF4qa7qTE8Ifrf3OBjfL5tl/dUqTJHRorReSJ2F39j20bfmoUICUya6yYGV0
6TtqJKfgcGSyWpdlMv5tbS8iGnFeL0M2Kg/I/XfGPOV2JAJEXh8h51IGUXD1YQ8LD/MmFDsMwlkb
wnlolsO7MIUaZVREtUOlJJGgUk78Lq2BMGuAoZus/EwsuPrTs7rmNj4iUKmd5sefFhFT69QLcfk4
5E1Nd2l6x4DNwKXlyUlj23q6B/zPV/thdsgf2QO0YdL1RW6HF51yv149pOCBq2b7b41kEwws1AoO
Mnpf+5X+CICc/7OD/HHKprMcsZ+e70bK653M4lq8FAz8sp3udwhKINxsE3bcn4eNczqYHoMHeO7O
8LArEm6byc9Ws1Qq4M9YDE2gWwHSau/pZA6f1I6nGQ/2EcarBE8n+VP5U8PtbU3/RbVNf04obeB8
x0fimr8v+l6djDU8KE8Sw9Ko4982CIIyex95fpxJfhTSyEL7uJi2JI0JvAYuf9guDQsugUf8XYvz
uVt3BrJY9RLBbx8SPWoyjHnLUNhbfOJmlXvVBoSICGAoiIk83kyPCMugCBq8KYHnwObmu0gZRRDd
sQS54U9OFX2oHPp1yh7cCfl5jYU9KNvJ39xyJyfBsCT8Yd8Xu/O7UpnqB78x+9deU599pfoasTHC
Q1ep/06/0pLxtmXgK2k85nXSbwzDfxcQtTW6XWzJDstIgAClVv1+zp/s8wQe2yE7TBlMzItRJ7dt
AyodWLlEEISsGNcSwXoWsq28tAcbECa6btnElkUITACL5UGL5uRaZ31m1iyLXoPWKpg+bX6DVLeU
SlfpaBP8amYSO59IYNGPFtjzkvQoXl2Gxs+6Sed5yRPNNVUve6cEZHjZMmnLSC3aaOZPhJlFGG6G
E20ongzpcq8hQyXzd/C8+Pc/rmPHYjh3KFqom1byuXT+eON3jFn/PPh8HYQmrhN4MtaV6i97MyqL
er4PkP+G6507NDeZBrh7DxPE2Q+q1drPriaarU/OuSPQbC3aL2hb0U028Q7lkFmXyXjEjKZR7OO8
10nDZ62BUmZZ0zVH+FGPM6pczpptb+BQWp/vLMpaqfUZucV7EKdDQ6ibqA81AGTTMEKZrUPNL2C3
0jfhyPpLU8oawUT4H97lPOwLhU6p9OkWI+WrfQfegQ4PIM2+OnDOjcEVNhn7ih+m6oXYwiB/Nciu
1+7JdCaVfML6NEaRFNq9/KKNpI+7x9GeCuTCQuAWXKTne3xyw1aTeodrt+BpGfxGtT/F9ronB9uD
+8ND5/1HXojhskpQzCE+0xvavUc3qOwgUnA300HFZft/TYNxihNwGVJIJz8J9w6g/rrUQsCXj3j6
i4B0Q71KIjB6FPGyvA72KhNwGQP0JmGSpxKa0yS5Upk2umDEm1Il+vbc0fQfglp5ROo4W3kdPKPe
R20rbTpT40tslhfIWVdkGapdGRn0srGykei+wh5VoW6R+NYAfgV9Dw5MzwYu5zJ0y5LpZPbL5bOj
I29VVgpRH1iZKCvVj27SS97sDFjxNfS5C0eIVY7//f9IdW7Mudd6EtwLoabKYp6jRR0rn3Br18yW
nAbNn9lCwoMZt7aIqk2+BA3K+CzIxviWK6jjpW7JuV+avi4IOwciIbDRnII1TMlNNIFcnWxxMa+W
yEXa5QqTwIbdL9GZ8vxSXr1lL1Up1QY6ljG0k8PQgYqKeMX7iSLNfmjlW/OHzp+GL3rT8R9sXcR0
VpkeTaBhc5QN1uJUikpwJB6etMiiDVf2NuITUHSto8BwddaAvaPNTEywIAQHZZyDIRugSWINzi57
QnT6op8v+r7Zb0DccH2muf8jVmKMLeWWgVapMm9atIo0OIff7bIxkCDW7i5bTE3ylVQhQfjcFNA1
dNbckAkeHqaP3K53eeIhqUY8wJh/tK/Qy3vB9kvNDlM72VQZXPBlAJt+DjLjYF5xa+Oytlg8rtkb
xqO0lVZUs6WJrQXpLav8ucFsdyt+ZOetncP9G4lTU3g/IMYTPGggTbOFnWhG3n50qM82CTX62b5z
LQWIkfrJnqmP3vdhe/pNjCaDr+oOZElH4N9ajSn7FAsACYLbm5s4kbcFY0ldpiRes2qhw+Zh8fzt
IWcS023ouJIH56/QMTx8XgjgjOAZz65dN2o1YO+Qnmu1aYPBgK4GUDc2ZxL3VHnLEPNlebFrn8Xz
2JYDKNCMRKeiUGCDtyWIZQkSCl7TVRxXt1QWXQUdSlzO1X7oHo9yJP7T98Nf1ZY38ux+L8RXnAbF
oaqSolI0nMUAYHbTiKaC1MucWd9P4jEIXBHXY+NyVOzVSx8AzHm0GFc+JyXHkp27dQslLVG0zy3A
02F9XBxB7L11TnGipeUpXAMNI1aOnJj6bzCmLH5ch75Qb5FB6CLH1uRLbaM3vLoXVL/10fPYWbsH
9BJhELtj631sqVAo2mTB+eNHNEfVjINE00lKeSMfn0oO8DmrD/nRBA/UEfi2YRu1Ex5LU4WYuETZ
mrfxl5l6hETmhUm5h4+v8tMmvEuan5bOwN+7dah0Bx1gTOL5fBx65R1VZm/V0wne+zYTnNOEgl2e
GHl4T5LwhrclmY7SALYz7QNNTihc6RhhCfobs7761StPthxDsP+LKcJewHEyaCVSJli9HK/xP7mP
tYm1v2ITwnkYBzE5OIg7WLbhXV+2IwmnIFpwaoFKg3LtuhMOcEP/fcpmzyw2vYjJW1d1H5gS06au
Vm1BSoPlp4nqcMYcU0/3SVLr6CRX4XWFzNQvbRYmVyoMKHl+BQPQHBs4OyM0jQ3wsFGDK/B4OSbo
duwCCCf7o7+vCt6pgkVQoSNntxqErUc+8YFAbiB4wKtKDYe4nFVFhTFDqKE0OOW31p1y7mL1UgLU
3sUeKVhvnYPh1hffBLGRbrrqT7eCEgYxgGTfcxY8N81X9L0//rTfTh0bYEMPpUCZ89D6nHk82SnJ
LdNIBe3l9+LrDoUWfbY/PCEfZDLqmfjN93nGVnEGjpD/K7PTUC9IfCxC+RsPco9jA8A7cz/5fcWM
zDB5bq9V2midrxaiWVLNfIaMhfzamqddGV56b+lNF5CnMhXtAaQtWW2UKCM+t2wrTXWLNtIrgIeE
NX1tkUKSe7414grYHx0zluIkmWo5adYG9HonrUYJjrtcOV3AHq8r9ozWBw3eVZn4Dx+x6SMBHiGm
jn3J+YMq0YwCDCWvIEFI4bkWWNTVkiB+qK7cfc/qprqUeCau2Kp+iOSADRg9UU6JLNlPZW9lgtgU
eVnkSB787E83p+0fDT5wUc+t74iSmOUw/1jk0thv8Slx7x4K3r/0ifoqXJvkAyXm8mozVU+2Rj8B
TJSSASA3/B+stLf2j0dS/JwE6kqdZW4VsYcVYequ6sYtxGfVryfHtaAjxQdO41OIO/qF1W6i12OK
94405WqI+IdkHgYyOqBve65vMXpSG8RphJIT+gLI9gIDb6h4gPucD+xZSgpDmliNjtLhSaYC2sCC
WpNL8bmx902UYaQ/W1YoHdVZ4LSyIqDZxemj/VPy0ktHTFALpmKRV/3HRqcqNkUR1wYdcHk0w0cc
+p+1no/nGhefLsDLzALthnnc0wOpKUbYxTxXl1B0nCE+Q1Y5rYNkYykwlaeTOm/O3wQ311GoLJu+
fejQCeSz+sTwiUw7jiKU3dboIoRityN5VuzR1LyZtCkduX4tsCrRDMid226+RQy7AkHszHG2DIWv
wBmgt/ReDiNK0/dS2gvxBSZX4yu8eQDLEjQhlvAgq0BtwKw2kDPacqIkT773pGP0R2oj9YK2rhgU
P3N6tnQSKuFh0RyNuVKGiXxICMacuh2Pe0x7RTE4SPoKmT4iH3amRKsTzBHUF2BSO/vlLYenVbbY
fGX3PqYURupvehIjvdbJhzeco5P+Mtz8pNjgyLE3Om522yyf0sTmKTnniqMfNF/Afi5MOo6TdbqO
k9rqSYfMr/2ssjbRHVP6RKp3wdnIVaYOQgFxv02ClF5ZG7O83YFMo/t+3WJDIGPpSElexMFo/gb4
4EMZX5dG8IpW/JCjxoiocO2Z4/kgpsIfpVNjRlrP9Xxo16c0i8BvHu5Y8Bwr20hWOgDKzOcEnecD
A2QFOhZtQUZEp3dgkzPOChBIs8TtKLm6A/KJyni5wkIhdKABB7pvCJ2bt4lpVsxRBxWCfoHehwmN
8VGYg/kjqCMYJGtzIGIBiyAX+MlTyiQ61wVAh8bosrwXCF4xMc+/L1eUX7Bl0c7MygY+4uP/mXDj
UZzW8ZJQE0WYr6oP1JPRXRMloIkyTEq85Vrg6x+PycdGWxo6DM9jd0pw5aq/LtpJKibLgxSvkdB4
Yco9Fs8eqy1nklnbAmlEGh9yulc8Ac0MUbU2NQAAwNXjDCXa6qIf8rrnC1q12T5kQzUy2v8WlzJN
c0QbMfsncu1f/Z6V6YBtOtLebcxVBm+ygRxawdOPhN/dWi/4KdwW9ZUUfQdoHxsXHXAbtEt0oU7p
5QRZpE1Z3KavyuU1KYWE4eDnAaTlp2zb8xifv9W9tTMLrwoSJZXR2qFVAtirLxmR9NXFRBztwyui
p/MyPjecuRpX4Gd46gxWZpEXMrkTlE1M387ZFOjxIK/tk475gFMvxOwZR3Wpy8vfEiQSQ5ryRP49
pKsqzm19lpB8U4QdCphuDTTHBWV/U09KbxjHpxa7qYiLxX7LTun+wo20P/nyNxfO1xuMN7nNdtL5
y/5uEcDMjiPfKAT+Av4cr4jNqoZ/e2HoVlrxUiusJk88H6Sc3ZPP8rfWHHZUzhs+yvZozfZ54X9z
l9DiP6K24jcKYQv0h0jboEhlYjT2l5nXE0A3gkhD5Nic/ch2qpz6MVFmVl1SnZCbNUcLIVDRy/re
NfV/36WZAiioaEKOqSSor/sCMcIqsgg46A3copJKjqQbey6bqFZORKdIP9Ol4jxJq+CtoZtGWtDq
4WxJPrcCAl3YfC8Y0QVJIWF1WLl6KnuaIqTzrPCF0iIw74XNwRpdFvlyguWFR8s+GymG9YBTiAf7
IQhy+7a0nyBk87x8r4NpYz/++bPEfgw8NPMl9I04ZLgI5Hf4maaUHmk35Um8Yc3wVrmbhzXWt+NP
hJiBv9siGR4n0DM8JpZeYNJ4a3uHcufXYj7KYp6Ne/sdrAzJnDp7Zf4aAIcP7mQYsvZUHlXPwCqB
RUdG05pvC0QOutPs7f7NITncSvrAPGVAgotm/igDnqtrNwWKOHz1Q/KNH75w95AQXeAQ7oVqNLdP
a5QJ81Cxzxej6k5ahzsfQKGsVR96ducBVX/xPsAJo7uKoSy49WMfeSHzeCfCCV0mO/YTRnOYDZlm
iH7uKVedw7MQjRVnrytW2qqVYFjwMfvB0wd0I+5Iw/m+3yarOJFdB7bPSLe2GtdCVUwYB8iTdpeg
4XHs9s0XeoNxucmtmY6tI2Eadtz5Y4lScIX0mV05BIWUaErKYKNf3QMTP/NtDZiESKFgbFWySgJA
OXfAWS+GT5uAfH2LwrOWcVMiHaMdgIyCdcCt1VjwGbyxQCWE9MJvdSQ0s+VU7zFiqO/OsSQJiRj5
17zjde1Hmg/blJS5OnJpNmcByw/a/1AxLr+zwQbKdNCjBeUWRGK37T5W11NviZDTzV++YFyY6hn5
4N+12HsyJ0YJhblE91OlJKxjWs0TkFKbd8Ar450vKQkcClJVR9SAvIvWx5fcTQzkj8rNxYiXrvzm
mUiP8McM3NLPUYz1EG1oIMrccrlxyk+BlsLiifi4B4ut1IdHmwXeql3TzimgHSADaC2pIZxGdVQV
7qwNt6nvnDqtRDgz3WXB46FdNVD9eLcXSEFbNltOQF4CXW6aLKz3YvJ8bikwV+VBngwCtAuH9skv
OJCUt/LcJFspPY4iU/HdPBW7Ji9IHpy7z0x5krqtY0jApEZN6T1KmwKqGb+zcvLzO+5iqqIPEf2N
MuP74aXSphpoqZ+iQnRrJHhobTrP7JfiS/eDV08xtkuaqldGsPItPgt5urPRmOcwQ+5jzNvvRVa6
2Sxeq7/IfGIdxVNPGYQPtIO/M24ENLPCJxo2aoAElrUaOKoVm/T97QLsFd9c88pMZgKBtBhL5XPN
0/Jgml8fCyIr1DsL39oSEi/svsbOHfw3aqiwsMes6dtDQhbGOBRlSPCjL9eSg276c5/dbIrypEwm
f8hwDQm5SyWFrlfzmloNMVg/KyRt5/P8fe896oQS3Xc5m302RnKXyyc4gDk+V0rJPoX/5XbCrabc
nop89qEY9zLcQ1HGy7MCM12sbXNkfG2WkGptgN/MUIouTooSQtJ72c08Dt+uyfBqOqG6q0c8NLi1
U6CMfntXhZ2FDgHbRqD4eX4+XEgHWE04BY6aJ9/h7JvBqbyNLJge6evnhe7K3XVrI4MWbZChhQK0
kPNa2l5DEQQejhqUu0kHNmBbJ6YXdKuOQdhB1PylDYpsEK0LrlcMdGAj2qChASkpaJjILUgF8vKD
P8glrFohArlMR5gPqbV7P5ltSmz5+74tvp9aqnklBC5ttqITk9Ci7X86qqf+y+AfvHVJSt4zGRZN
nGl6G2DUkK3IxGggm5rtRurw2sLDnqNTUnFzcfn7+OMT+zTkuko68taqiUeUQIEwbMwWr8vHKevh
oRgncWkEUVXvpW+WpyaQoNVEfmOTECEakRNQDMEzIHgzt6N9LofZZemCQ1IVsL4PfDltSbma6XNd
ZgB9eL30YT9s7jO3Mlqfu0l7LOHyUwU5jBhxpWnG/9vQi57t/AypTLn59YJFDA0wjnb7R48BkEMH
aRwP6DJ91li5Uj19bdJL67iEzpRwAjSW+35nJD9HT0Yq3I8V1wl7WvJtIufyBERbPlvUXxuZrBNW
rIzvM0onp0dz/EYl1bXrEP6fE4RYiya832hjlVHYDVAxJlc7+npT+a4bkGagodw/YstNmp298MR8
eV6vSalEs1eiwB/43gc6ralek1J6hgsZA3n4El68fszi/7vXdWl+Ef4781ZAjekK/7Pycod4xqO3
2Du9FIs0FK/n470WmeKIuJtl9OsjeK31q+BooVWpuCZf3sVCR7Zgg0Zms2n74UITbAoUPrZ0ZaH8
VYjOR/ci7WZEsp5Vm4nwxdcVNj2cBPbxpp3LaVsRj79cQzZ0g3i1g9aBHnDexTqDR27KImlYBOrt
RqA8U9BeKlarift0jDZ4HxL+2fjLSyu92sIAn5cXS31l3wpbuFwSDIRahE9/zv69dGfV5lA370PC
PrmVWnJCnm/+iI6Rw6QKuU4xAFWDNVdHqIqSIsOFlvDYYX6oNannJhK5sL8LTdjMIQlFXMHJEuwi
T82hHBy7QisoP2VWH0vOO/n+GXLHxCxWqDrM5G3+lNiR1cRC+EOdJh2yKSf5f1/SxBtcNsQm47YY
VCGKMowsyLBZzG9pD9fsyxYfWuoldYPUV2QndPPjXUKJrutI2x+EGbBi8N9biod2KbHR5q1WJbcZ
G/myoQ9K3MMtKMrL5VLWOh4aLAOCa3pRm2v0aFi7xOtftCqxXwT/AvjPFxhPfjN/Ku52Q/HrFs6p
pyM8Z6ikSdPmIw3VBiWH0ExDF0jsQWdKc6yuU2xlNwK8JEQYuoNpfBfIYU813Pyj3eVLs5+olYj8
lMHcRgTp1q+ogou26Q85JOBcdxjjMWrGLNMHU0MD6JfJ/KuOeg+F9zLfaGYwwMwPJxuN9NQjJQif
qqAKqsAz4Bk48GKB38CtqouUDr1ttZwL2amCEo28+VN/cNLhEo9TJJW5FMZRe+2Q90ziCxTCEP/z
TUwcNop8SeppH/oswMgfV4TUDUqpc/TAT39t3BHp3DLzo6Vy95jQh33UbEeFQAi3t6ZwRpTZQvFF
bf/7XT70XcVgcLoy0UghQIA0l8SbSxFU7IkcrGiAcWV3rpzmK5YR+Ylpt1eQzc330MdLuO2NSZu5
QsYrvh8dK+h5O2ACWzsFeJI1KoeCdDi3JkgKsURr3QMb3kw2MbrND0Ydud9wjQCrAyfuoFeJO/fw
+2Rffd0srAJQ1czS7QmvhKx9fMYe8jEw0CA496VG7XJzjV+7IZic59KZZlK5BiVHvXuIVbr7I48F
fcsYOcEDX+zYYvz7dZ9x2KatnHugogck9i0zlzHyC8eKgich3rCAOPkM+TUBS48Y2uMHjikhYKhi
8WPazBh+JQV2XRXcDWZveNCIVNIpg8wJMc2+QCOYNcRqCdfs+5igXL2cswwbHtZebCneAlDqfmIb
4UtMZmz2sxhREGhKLzJUaxNau4mhzEah37IkldXiP86v2+z4d86J79ZrgwCDT3XSDxmpjJ4Q7BDs
Uj/GcEHhkRv2177nNUn7nu3EG59keFQZvjyyzDRAL8HTo5htyKB9Op1smD0uTv0LWilVM2ZbfAGi
RWLpIS++nt2TkjQqiCQXMHJ5ISvITIenfUJ/cm9ScGx5JXGP9yHy+85WM+rYN/Y5iCMgQlC3vCEv
XSOSCYCNdJ8y9j7BDbotgoPt0zj+sW2Ena4OBv39qYxP+Domn50G2fO1qxB+hpcjk7rwexXfKudd
6WCoQ194ST3UzwMWSYzC+7NB6ri+mN5mNJUHpHeH2wiofoCQ59GHmCTHrKqRQF1g0UyFNPLIO0ZK
uICKFUid28vK5xymbQ+avgwgKCXLdlzOW56BeY5eiI81y94U3T+4Y+CZ/sEKQPr9DU0mfyelvz6R
7Djo7RbImPHYf1jbBVuNOrr/fVTozZhadnSDxgcjvCF6LzUViEhKghCB5iexoKkgfTCSjfH4n2XA
/vc9gsa7PWwfc7t22NDzaXU9Jc0Cb5HdsEZGIMs9oiIdpwbW8eqrWilU2AYkwbcSwDwZVHfHrnZQ
Fl8tUy19HCjJP6d1Besk6W51zoXm38FuIy8DboLH79UZOvaEWI3A1QVYkxdlSqJXykkFhkytWkZk
905U6JOR+RI8g+FNswFr1sB+W3s4YazeGsoxzfoShgfZdnc7SLqB7snPQQmcfyjnZ9HoZrxrq5AF
Sm7b4+6vi6O+asbpXBtvccNhiduNf3jITnz3uSOTXUndaf4FpXgS0qDTllXt50aR9UTTsKV4W2Ud
/S+4F3DMTC3TU9eraxjlAw6Ttvu8WF1MewExJ2s43wUYSyq/je6/FFpkot2mPRUoTij2uoE6qk5g
7OteKWsAXpJLBNNJD6j94PLLkm/62JhIDF0o27tgtwhGZZDBeB2R1/SSWqyMLrC4eo8tMKS/Iito
L8JEWSNvZIVYP6SsHve9HqCt23o63jcF8dFow93QKKFVFCi1+FTodxXTRSHlyMcSHfeqkMwZLl5h
SR1MKQvpYRTcUjcw+7aLztNCn81PtAhawmscesiUC2vLOzrVuyQv6euwVWSoS2nhnMpwMTKyWf+x
clDM2Kw5bOinjyQ3Z6xTRvL72JxquZ5EOaboDSGNDcWJ2d8tLdVDsptiMzw1TO5Avhg6RTR5U+y5
NObXPhbMA1lDsHUsecxx31+R1cIPHt9gRvVsnIxhOgmbwiQtY0f0ZJr9nS2kJmA2zmCzBbXUewB2
8wyQ+DtrU1IJP+Jch7g/ZaE9JjxdM+ZIrXMP85h22uH2pr53dUrnEFzR8B23QOF1joJQALEz6bY3
0Jv+MDNxgqPGCOIO1LJhfZWISoPURw09nEcWpGnmPzOmqwBk62Ed9CzmIm4ji6YqhzZ2ZF85LZWy
9XcVnHfB8JKXIvD3um4UYDskJlbiwsm5086Dy82I4oBEJXo8JOhzIPpStNiEX8/IfpafCn7fnSHt
S4jFNg1phEOmRXcafiHwKlOtFcbOXbcyWjinX6dxcsNSBVT9kxqptz47DcQReceVtVmiLjep1qX5
9yfg8f71GmlkWoOwH1oO8RfBiMNqUMfGX9860xJTIzk5Vl21KWhZJiF8+vDhQJ71HBr/7C1/h5tX
7Q3JZFz7i3KzDnqxsiUFrfl4twc897DBwOE2ao47FhK3wZzB2XBd54McHsHFKC7spzrlUBV5nK/h
cwe3ROtPHQ2zhumhxJ/qfhKs81JWHqyxMSwjnXmScHCyKium6xUZi3pual6CRHC91YMkYNsgncxZ
QbxRv0VIcO5kJrdKehU4ixk10QawPPtNgTLO9IvS6Ds/lF0Q8U6bV46b8VoBLJkm1uD1hHYRKUV+
Ep1yXVA/8FiWZGD9UqdrEnpfE2iLdtQt/jBnMqHkWEgY9vYsHmdHnRvpKpRPIFuhA8OaTpmtgFC2
I6Vk2+vGaRKiPv3kErRdxIVf4789Ublde0adQx9Duft7gvZwuwpgDxxpE1EloCSXE/bgiPFqHMmc
nTbazb5+wZo1TVDJoaSv2G/5IIdTXloSM3mVzERB/TnoVnpjC6bTgGrNJ0x0SNFKd0kf/XGN8od5
VbaQ4JxGaMc8wgI3ZMESVfVuItFbG3AqbBv3T0jTz0m3GP49JYg6jZuIixyVd1LmzBMNjK0aH9dv
9/LttxPPjlwfvIZp+fqIzkvMM4fFYMtfAmNQ8poJ90wwBX2BGSUDq+defBn31V60r4IDa7DJ2hRJ
w3qtSnG/n5lCSPwcnxiDIfOwjUMC4fEE0mOom1Hms+Y4Jv+cBGn5LMDbDl28pElraS/P7KIvmzKt
YDA9m2QTVVReLngGNOLaIaXXKohy5AhjRPmai6kE9Na8LEIvsEoeK2isoiYrFEdUeTzDCmFzmYaE
rXeB/VO4HrZg1DOld85kN6ebhGEFIMSkLvBiRqoxZG947+HmFWu2BBeq/OAGg7VtjZ/fokUKILy3
ln4MAbFMSJrEJFV71h+2oj9klrWvqpca45UKeU5caorRBHc4tLmCH6DdIGCwUUNWxX9bhnS4tr1h
yzDY04+fk2pA/FlI62sx50BKD46D5z1CLDHg9jbMEo/oAo4djKfJ/YCuKgn+NGJiFJlsds+FxD8a
byJCHg5/uuJr41N8xn0XmRj5D5t3c+frhdWzuEq+ikG6TRKQcN3ErUuOwkLeg4GULWbJLePsvBaZ
RoTLP2vXNDkN3j6cnyuu2Z4XOpMTakZfg4Fe/XctwDpFty64XAyofN6vIUuqonxiLFb7w/MoOsrn
Ge+aYXsWymMnvfhHSqlFICLyJNXXVIeAnmsURPaWqVyXYyKjDIdKn0zoHEAdbhY52bzslDkTapww
8U/4tIyivL/FtogJkM6HnJxuzvtcEHbq+SRoFssBH6/xLLg+9mw+ljxw+u0Wy7y95Rw/4IhtU5f4
/VpzC0FTz74hp2O+UuhFKVcd3cczRB0VzjheZTGYl1y4bVy9LAmem09ebl2BeIq7ioEkxDXMTm8N
b9nqYH6LNCf4Iobrw4XuR/xVgdHH4kaZNfVshnwxtTALmQ4aOHBO53Ex6UBicnTF//i+jXzBrlZD
DRqZ9/fIyw3c05dqrQNBBI/El0OcuEYnQyy/qE0ISFVqItbzXXX2SKP6DBwB3H4NksxnWcAbWqGV
g0Uq7Jdyb5CuRp7xTx8vCbmNF6sZFVm0P/YMR+YYS5s4hN4ACTXfa0xoej1GBbX8zzA/BznQmgIJ
MwMd4SzJaD9h+IEpDsSd4b597ydeIKRqxdvAzgAjiNv844dYGylJHyBYrCcl0m3n0/ht8gwORAFS
FDURwARBd9NIbv5j3mZOh2bR1mZDTiE/oLqbBG7u7CvzA2enMRUr6Ju8uxxzWeMN/ulMdHoP7UA+
dTP0fQWYYbMtTPZlWMgczw9l+SXPdgCZ+7de4OVOs+rJaHsmvs9Ii/ZtIgbyr6/Bgx4S6v+UUoWw
1catBADfVwmH4BQcOmlH+wAuRWmWy/Opuu2/Q22yJc7yGYkeKREA9zmgnoaarFbCR3UKoUlFxm/L
GQ6E4S15d3gNG2qN8VrPxt5b5YFZv36U4fQxvlEfVlWeCtOqnfwvc8V0VNdblmcshLYCEf8kx+4v
Gfi6I7G1/Iia7r2E+a2xIiy4PWzhxwDsexT4/OyVjdzoKCPnEuM8xKqh5Hs8qJDlLdK4UtnViVGs
Nc492XYwMsM+0ijlKUsT8gv/bPd0ggfpjjNwhaX7NPjDxKZJ6EB8k15ETkrNVdxQuA7q5Fde9qw5
jxpg45DeXVWlTqL1rCQ8TCaMoA6usO36mwbVT5biksrK34ZxnUFribPgAbFYt6SfQrer7TTYi0jF
6TkhjlLIuJK3l8wAUtvWAt1H8bu/0LFXKRR5e1zSuyKMjbSZ1VLwls5QzGUUhO+pchzseYNQYQUD
mi+7IUy5ukDzfyMzgmcvmGTywk+CQlpUxJ0e2ylOA4eoEyu8AoY6ID8qZtKZgfzAdsl5AHSM2uop
2y7qrQUfPxd0r9G6hxCeaMFpEfJaTzMxJ/0uzE+zjJOIXy/ojyd+zdlyQ9+xRuraHZGxEsWOtw2M
paF7eC78i/7VWsR0zgXjj0w7kLW84tOglEZkSeOSadZeg7bMOpF684o4cFl/qbwS0KiLskhCDtFO
gJwzMNVfg/fWeBwpOLFTRNNr09OINC3kQwP0BWxy8cuboj5PWss4ac2rdB3f0SwK6K+HNfcAd+AR
hOK2GyJMtwIlvVxSrGDZ2+SOb8kOCU7pjicujVz+9+14kOvcqZIzsj90c2Pd/enLBGYah0Uurm1G
fP1Dd65AgFiUokA71W1EGa5zrNtQ/fD1913UxBnWGKDVfVD0f+0ITAzOdMEhJ9zhKLceElYYiowV
YbnfrlwYTtuKqD92DAV1IlNcCb7FmIG5iiGEUOxHf5F816iFCMJo1Vj0EncYSoTZTzf1Wlgq8FuZ
mRrEBeztPvWW1qYtQcU+lAiQ1LrLJ5xttakRAgirBBFZzIBAV2FdQ/4UChOdymbA6DjlKzV1QcYY
PSu1Mw5jTxgMDxldqqYGLVlM8E2tL/J3JrSHXeiNQcFlT6pu+lzWM0t99M0KgnLgjyQse+HUWex0
MTb0cFSFX4kS6wzAjPYCGPrJxZHwYkqsdruFByfZ5bzGsfWJOSNHRXdf4knlDsrigZyADxYmST5a
secE3TcSKxQnhfFX8QXoeF1hkMUpsg9XpoqsTV6K8euz2B1cZMppIAaP2/C+yQH77u/1cZkVVO7u
SIwUuMOd0tjBQwnq0PsWjOXjEQ8zetwJZnJbP5z4DJZ6nurWiaD3wyzzIYcdd5c1/Q2bnzDzdI2I
6yBaJ+AF29VVZEEiGfVR9+riwGy46MMYq2enIPEI8kQhZXeO63bix59D5M0zWK3ypyvx6nsbUENO
go0Brfw9CSq/kum7ySODTxKhbgUDbcMfPo7VP8Dw5cEOaHpz6qeYYL6l4dSdPka6eF2VmEPwZ6zj
BSXyRkjYcuB26Bupi1HV8Do56zMAgtumJ8lvFjl8TTkuMnjQKEyMnpdU325lCwPtqSTajttktRIC
6YmRuOjpWKaRIEDk9sLQQ07eKzl8xhO35jBxgbHPXNi7B7AC3WKrwAeSfcBwHpZXw2xT5T6cY8O0
/myP8jRH5pcJG2gO5DQ173cu7SiQIj3YQSQqSPr+lgijJ8xOo4fzkDlON4/3sCefXJayPZ7X6hXK
MJEqfhAxDVy1JYVAiDK/sFxYzwmHu7vPjaMGyd/sd3YlmjHZYDtNsS8U+fQoSm2lVdGCnER/8dN/
X57znG/4BVFNQ9aRWaMZwWFzIyr+SG7IiKk+IDW8PVnDjjo5hiimHSQ3uxADSUzG5u8O7w9z1D3C
XfUc3mtsijoKJB+Y369VAPAER7uBW/G5YGUxptp41moqOkK3dbxTDJYCVHSywoYEjJKHDfVtIUIB
43GwxWYnwXPJCoUeY1wI8RKbiMh+4ekCQr7E1PeqzBkC7szCC2n91l4+LdAP2qMw2F7YsZy4zPwe
er1cCb6DjbsVaC7zzutyWCNWznTiH4HbpTLa5BV790wD3TnTFixaX4BhyATwzL5j487XWg/Es28d
3IBMEMuR1VRLb1Hcl2zmH+B5TRxJ0knZjbvzs0TsuBMk9aZTOJbvqoXS1xsIKBoxBUnrFEXx2kUI
dWl1SSihnD55mIJ1thGVKatg208tFatUgDMoj/In8Q9YFm/1MpGQBGgBtR5PTR5VZkXMR89d4/U2
Lp0ewiLS1lGeOBjpcOUyFDWQj0rBJ+x8cqTfP7yfbNSFb5nBQT7R8TmhRSSphLBO/1jZLhssUIqa
c2jm2vB9F40NUuyCZkCtN9lUNHC/jr+QiP1Gehr+IIqJBY4Aj0lbguMTmE98zm7GNDAXBy1d1Wwj
gVLYWXs+1HSzy2JUzF+kqyiUEE+Hythn0N3ug4mLvSkgcvfy8bJTM/756yup0aK4hHKKpD4ozxu1
NgzRacyp7fZ9TwnJ40xYezjsJ2kOS9kzU6ugS60YV1CjafvK+h1qqrqJ6dF9hei2jHaTaNW0/9yZ
4ySX5hRihvWBsxWqS8jfYsWOpWnF0k463Sxu1iHRIpLHpFAWOcccDn6aQh5RfHywAiicsu078Ufa
qW3LwQk5krnR7vV6e7Aqin8mCBKIW7SMQn5sXSdRJEmt0wHhG8oAjeJ10QW7sKvZ/D1KgX0dn4yb
ABv4dlGbbAgMimtTM5CKk9V9tALUsQUHFuTgYx3L50p4uzSObiI24VZaye3EHpc3ES+ueTOx6NgI
7n7jRNRp0isRL7oevTasyGhQZCQqUFm3sOW0BZHPxN4SNZPJU+sAtYYBieIpCRAQGCHybLDf3aUB
JX2B8Vodiei41R7Ohw8ocz/YZ5wojgonzUbH08YUrzDeJDAHIGdru12ynYAvyC18TtfLWrgPh/CZ
dPsrADkGsX7dLE6/hEwOQO14MIgrZCVK8arUNSDN/QxC2/AoMRfdJov5kcoxH6CXf2OBT6ApIbtC
E0DgARkZ9mBkrHLyx9xIorC4xcUbpLPM5hU3xhmQmk+kMVWgfngGBCPcS0eh2D+KXeDETirE8Ptp
PjishV/3SK8IhkM3eCYheOZaiXa3gS6Ab+G9qTeQztXZP4Ti6H8yCyXwuI8AU+9WIebCk1ZClji8
zkhfEtMonXR0+gzCJBGiuQq+YuPXRMu6cQx+GV6Xu/tEiYIxlJEY5g5jR6V5kN4g10ObCHaY1+RR
jeMKbaCWALWBzNbzwpcoxfPzFKlY8HZPgeu5g0NutGro1VS5BO75JVfC4I4tsF4Rn+ZW2WmhzLCJ
TRO/FEMNcnywU/rvYyZzYio6/YWguTjYMFIsKMc/MQw2X2oxMzUqaDkPM0V9UgHnM9wOSxRhZOTx
XzMggLKJYJjD6kTLgnR1hG//Ed/otGqnoqviCw5mIvZrAZ+i5RmKizeWEp9gEzwDYEOZaZRuyI2u
LXuT5yDTIbDIvCNTXUfBzG9iIRumMY70EPrAQhb/HYAe/562Ow/DkaoqvPA6iTjWqAA5dSTuw0E1
i65fP354ggDT1dTaaKeJRyMmVWWoa9J1MvajbP6UHGQ4BBFmAcSN2lIzgE//RkIByAI+1FVoTrjv
nYkg6rHRIfRB4s1qZMlkPpvidcNyksvTT//wmr9IhgjwlJ/+TO8rTTAw2zNqD7dgNS8o3i6sGLGh
/KM2ttLlApJKIxWLRElE5fvLvcWogC/mOlduUBpHrlwsGBKlep2GF/Hksk4xt0bMy8rANBt22WbX
BVGOnuG1Cgo+GLgmayfLJp3wU/bh50AoZCLAG4lY2NEX6RmtvpbBP+1vPA3ev5mWJjcoGVqMMyKv
U+JcnlUqjRT6jr3+fFkeD0XdbOqx+qZiSh+fYfdA0ItdPB4JVE1I9qSlhv8WTENv2MIB3YX55ng2
W2C5VWE0+rLSKrwwXFugc77cjx4xb4zZ5QjxMQ3CGNa/EMcgDjioEYql6HzlJ6L6Zw4ratk3oxVF
atrV8mhK0v9cFpZW5yhrD7tazb/TQzSqvlqVxdFbr7uN939vkFm9kWGi7flYb9txK50dQmkHvBPR
vYvR/dbwYqIVzUOH81Lc7JI+cbSRhH4qeGyo4b+l4CIYw8N3fSFlEPlJ16im1+U9Wc5/5SJynr78
cDAbwIyDnOTXWfvcxrU0C76R05achNMo4uH5vkdzhs6c1MKDj5Qd/HI1wU/dRlrhwyZtc717Mzsy
Vjm/ztl3tt2d+ws7sGaDrzLeE2Peu7ylELeotUpIM+vldS1ukFZCfJ/ne+rS79twIvrTF/wL1C3Z
jO5g0BDzGJDmZk5t5UXWvIPq+5Ah/S0rq2eCoF7iCgjnYbz22v+Cequ/wjVOKXauN/NccV+EXjBN
DIjj19gy2jRi/hySbIpY6GjVdnRcML1/qrqcNDdo++2vAT7TKK0gZzoDtiR+fWxMii6pNM7cWGWB
HAlPijgg7afRm0ekvViY+qdzS2GILBQZmFOQVb+WS6TfcyMKWdBaeU5pIN1GNUi4nbYqkd5efwTJ
iBn8vgkpI2o2hVVEOuvo+z92zy1f63/iRPRxfWjY4/unEIKw0zGEGpALscifquARAGfv9AXO/TjR
K5kK+nVb9oz5/WJH+VvDI33SNignSFHWWH/R6ALSXX0O8bWnjPoS+FVlM3624DWN72UIJumNo3A1
J2p75k7EZUV9iXoZYYhXUAbhDwcdze3ZdgE5LZoyY1NZiR35pWHs+kx9UYi7twd5XS9XRXvMBzUZ
FIZJ9a+jqh5KqrpsZhsERJuSz+u3TbBvyJKsfv5hEXQiTCISQzWJACAEt5OJiE+0fr1P/Mqfe+wC
Bn0c4R+JnrLVKe1KHzYYoS+vEkaikdnbTgT6hBZzyRqajb66ma0MU1PN61+PjNS+ECgVjdLtJHp1
I6mANWuWydT5DIbWprVFCQ/ZUTfPpA/RxReuNmlRiEwXSKFX3VCTc3KiApRTVTe/ehjRfZRNmLYh
rXzSoRLkntKC4lYkrg2BMpkNgb2DwwYc7/kysdIF2KeGx0roqPuY+zQNQL6jDRcTDLZoBkei+OWr
JSnL2ShP194XSRRrSRxBXX4sonqbCWi/DOwScDlkBq+qhe56bnyVIHX93y/5Q7U/k/m1uB9ntaVQ
JA3PmratgPXSjPz7aWbAG1OVfs9YJcfkE2iRSsSDwYSrCCSlx3kGQANTKulmQndkizbcpAtCos8c
X0lrPC16GrnNJ78wBapGQdfRDRITuQFePjdzuzgz+8+VGeOa0YeDtdty2LAe8fhjQmq3JpzdgSMo
OK6EQpeucESJJT1ksM5HZhMCyRq/mq3i5cBbsbLK5XX0hdqK9hK1iTlYbU6fWzF+m9quoc9gEs4g
Cs1mOOpMXK79VcQLd95IcSZ49+E3phpm2vnUJj0D5prVOorgDNX6Oqe+ViL8TOXsW8snyfIWCh/5
wAElCD5Uc0V1CFtCOaRfehA9WLXXH36lTZvPjeb9+lxMcmortWda8LAa++BpYhDE3FZ1ifOCljS6
DcHATDFOCMjVXzXOaPzMQeps6ez0hrOxPeNKipsmoyosO5wtTXQvs+dFFGBnvaEoUYH35tSyh9EU
a4/1zb5g3rTEUKG+YfDMizm8vfTf46kTHdfyfK46B3kOqSvl6nqaxB/he21tDoIk1OgExrUPXrby
g9bmDn86qPV/FU7v4It4lWOoNuT3ss2dmxHaQTfHLH7/+7tRxF3VbxwU3KFFnouosXelcLUvoLkD
INsnYMveivnfXEmlJ0OZBscyexGT2szKTXxbu90SHbxzMay8m6uDBC8zeli8yC2fOd0BVzopzsKt
T6trILGMCIWSD3j/fahQ2xlpckW7VCnI9RJZNom0qB9OcOwSgFcb6me9h5dKUyBcfKgbAlnbZvF9
SDsweRC79TSnDnwdRBD18idWXnT9q2Tmcg1G4QJ8slzATdU+vISDAKowMvpTEEQ42araFQz24Mjl
q8SXkqA/OJrmb42PGhyV3fe50Vqqr3qXqUv4sGxcFtMAXLFjo6WVZxbZlXWYCoBdydeBOv395tyk
ixQYr9+oUAfDIr5TYqzYVbFg3SNzW2/P+fAD5mNHZAmmF7NOB79W9B4PNUH2p16+SFfQwQ60U7Qp
SIgXuvLsYHZNMkAYeLAMYdww3aRQEtT36DvxY3sG2Gu5wF507EdxaIxdYt377E3zZcfw7+toFxVI
K9eNfvxbzX3m3BSws10uQk9bVXZvHoFTfbSqgXJLbYqTtoloEoJ0qkde69OvQlO5zkWLSK1+2HNM
RuVZvmn/Ot+CQQfqc1kDfg9U3xuwFV+OdSX4mV5fW7kbihXosDK3ke0rh2nxaZ619iudLTqJVign
4DaVI49rp1M/jNeURdCNYw2rYrtiiKSaXIa0esy+UOzXMESRrDfg7oeNJY+mYxtXcYMPCekvtFYk
lh6s+QfQxvz3b2vOWN6gStmrzPtfr/ANX9G5sP5ldg4p01XpAzuas+cswel10TNZbGOdh+gHTQce
8QHouK6cM6JbXRDZes6wpexaKAb4H7OSuGyvt8MzYKFlMLry0wz5HDmIOdsVmooXYCufVD6bRcTw
kfl+Z+goz9TZr4/SaCc7LSpsgkY3M1vYW58KQQDMPD4sK7RuCuluymp0D5IIv8I1JgKFQQU07EtE
b9VfcMm8e5sC+Hro5X0m8/jv1vgWk4Fv6FApyAT2dK6u/ejMZ4RtBogy/VwBJ5AcoKgMZhkZJW5u
62XsRgksM9dl2jdOKrgysepfPyrklpP+qYg8SjqoaXImI3nrqdNvjY3MmJy/w+fMJJTB9dmC2to6
H5mI338Y3HWFqXE/kG6XQ6JvhwOo7KSr8SowXhvorQOc3H/Vkp68wwRGCi8U90Y7YEvg9SDoaaZo
d4lYfU/S7k9pwQCYNUabi8erncNoC+CUW8NSOD693SF9EpkVit865sKxmoP8M3v9HDUhxAwpFUx4
O3mg6cxfF2e08IrrNccJYRns/2YarlHa4FWtKzkvZuYnOW+69rjmNE/417REsjklf3Lh5rHk1hye
UbHY/nbIr2w66UGfCUPBT1bzLSGQQiJ6jE3PA/xYgbA+bni92sRykBLEknT2Y1hcb8gjyPZyGsVR
nrfi4jTNgQCVy4czfxcKJfOOPCdUYGmp4Jryagui8sSAm44PG2e0k0loqKKInYDt/fMOJkD18PwT
2dd8/zcmmL9mOA6vO4vd3S/lCPAOu9T+slUJPEmBNbTz+FnRN0MH52iElaT08JSYRxwDXbAfgULB
F8IqVo+Zpq9meH5Fa4yFrsgmeI4BsObF5pON8cnDsJO9bYNyTgmYCBXkSElD9BQyur7oRZs1VVd4
7nBoewIZENmId4n9UKg+qFCS7/XBoIvvzr7biEQ80AgzIjUeEeV64A4uP80dKiww4OKM7OWM1e7A
f1coEGTkzWuCDbfYtidndc+QIq/B58HzLO7V20VCt6e3nnRPg5SCDfkAznelIbUHq115avGVLMFA
NbxqLUOviLVoilOFQMYJpEKT704s5fx4ukPr+z1Gk1BfoDo9N4veie93Yc2P38yFTY3vmTEAUEhr
eNmV7nWyCUQ4l3PT4C2ibrJtUGh+3i/2EyGoMjGk9phpIDhtZGb2D/eFytMHpXDX6KqXMUEQKWIk
aeV/iV4dYL+HSZNnfvv+ql9rqS02epd2ggAptICa+ziL15Wt06pyp4PYzHkisC8IafJ1sWGH8Wjx
gjkF9nS28HR8YgvE23Z35EI8/kmcTqvClXEtTcD/SkTm+CKjA+/hGb4iIZmnmDHicuCukql6Ehe1
fuSk7drrNWej6hZ3dwTt52mWY++abxKhZ7dCdy3n1lJjwRSNpIh8FsTXp5fa8UhCXtlnzGWmvSb6
ToDrv4+g3GDtE1zfEViIMxLY7bRrrTroTQRFy00bLQvhkQmxzB695KgguCmu6ikrCXod0v6sDcQy
UPViYyEFoLlh1Zl3UigYV8tyv6diJY/r0HkPif7r7knwZXPkGMQD1/e6qU2Au+GZXsttuPrCvBdI
Ndehgz6FrbwNxnRlnei9YEr5K9XVnMIavLjvZ6ZAwJsJ/4jNgtV7flap1Ety85G1xJzPfbPHYEvT
G++gNeESlG5b7rdcVSGNP3o2pr63NNd23I6yPpyyjuLeA/7J673q0P7GkZ6iGIJjC5olMXWd8AGf
YFLIOvpAIXW6whhtyJjUS6Q6SKimnUZU97h0b+4D10zw6WIKvOQH7KfWG8xebl1eAx7hpxaIFRVe
m9YdHB+UHqAU4UlZI2MYhK+o1eGPvHdVq5V64xkkIc15K1D/XoiQhk6pi2rQEuXg/J+03KfBE07+
yth75ByvWBGDdOnWY9cesTwKEU/33sHA59fxUfESarH/bbpYGGsy9eifPoNMG/c4ZjyXhGZQHTBM
eQHYBKyJvwmEbH6gdkv/jzGDVbKhUzBvPFtPcTfseKP5HNAYGPokaZRP2zWf4sLpwlqZubymqS38
OwAwTBZ12pppJONMQ2H3heMkD/EG6+dvlirttbfQPrJrr0y7QSPWsfvaoCcjp7zzOyAgE+iVXS4O
J14BpM1a8b/+vw2G8uUkSoYFwKuI8BiPk+1FmghcAUOnQqgYbV4kQbXJzv42Ycr9/obB3eQ4t4Qi
WP8g+vrR4OL5k+iJ0v5OEFTshIDPtwYv8rUKv7ABwDg9E3UfFuW00y7w2hAjSGslBmNvAZG6nBJL
BLKKe4jY5cq10Ze5RjmoBjM4yU0oc6EZsTmQ8y4HTpDk+e+uV8nAYDiMuBTqOOQDIWgn0Y/D8Sca
AOVUlpDzgrQFy2oP+oUA9Pfl/fbigkboRKXwRFbIp6kCvGKQbVCysachB+qsm0yrdhaortVrl0sQ
Mr/w7kBkJ/1hJuRSW84lCsGjtGZMvIYOJw2UicnWdcNc9QmcIerH/eQAB8+1xXyy+FuV0XsAtLZE
p8tlQdkCvpfGNeyvPmHRfcfVZQ6L66MzhyFSuzrDK323gDtuqgG5xjRMnqQq6qNn1P667IOMimoM
W4bK+KjdBDIKYzfivjLBfavJqQ5DmJK6279zTVzNQeg2pa2RlNht2DkloUc1Y5qpT0ZzABcvnXYu
0XzXqZsZFyYV20JbzN0+EuKoYAKoU/5tnCetmMY/nGAqJXlSe0fMHM9MuG6vfYFBAS4nOxi0faqe
vHpDFvus7lptuWkUqMwjlFNcGWf0i3uMcetVfi5kIdU6xh+xbCmwfVe3H/vj2R6o6Kzu1lwZpFer
dZeBjezmbzQVmaBJDxhfF3aK5jlptKAIrPxM1S1wBw+nzBO9cuyxWOfV1X/NMNoqHrnXd/SZqEPd
IfhR39/FA06O7Eai1cvw1NNQi28Im6Y3p2B54Cktu4CTW0A0rdwOzyLc35x3AhmI3LiIZNnPm/7r
ZzAaUz/2C1OKH/3P1ledmGSLeaMf0gauDDueMGddwofJBI5pzcagS13lnOhcESz3/5mfuvZfEWoG
479ACxD9w1juyuLRnU1V5E6917a1/vgb7bacGdTVxUy/kljKmMP0rwUL1uzGTiA3AjB8dCQu1qVd
SKu1VrKivbFrPJ6tFSlyJ3ShkHCoF6JIT2PF8UwYLFA8G9e/ggzdb1fLwhDoXeyhm7g1RGQBCNtv
jj7W6nw2a6+ipwOB2SwisAUE6Hzt2Fm7QMW+aNHuSUpwPfM6x0Fo2PYqO6TUZpfBqfd4BfPzdjPA
BgVDFVJnkSikMW0hojs0tJI5vdJfnkpWTmlbrX5Jvg9HcIaXJBASp/CTpqhwReYbx0aC6tAwetGb
Vt7XLy8k/pHpm4uRXGwT8Pbzby31SlxuwGprLBrRbXHryrS9rjLWNhZIyBwUT8fXCIOVZhzKSBnv
wTyCsV8evccHKrg5SggFLoQ2wiOxagQHcKe5EMfttLSwZ8fXpGQ8orCJ2wkDKztdAAHYPIKl6kAq
x0e4nQjnxUcSEyz0hJnxfDTbodK2wkOOdlUEV6ZsF56DjV98wkX/Rvv9cY2hV1MGQHRX/3jutkrG
R7F/V78k6w6qWhJ2v3On4UGjw04ycltmsuKrgiDVA2zneA27eTXQ4Rz//2CC/WnzOvpI3NXOD6yC
HweVdsTNjvIQ53erDNxAzKGzRqMX9iCKJJV/uRosTU6XA62cHx1mG/fU+JTy+cho13ZqjlHhsNth
HdWXY6tL7cQgJIfDhIvYUPYWtFVqBv1tSPTTRAF+/p3D1TVToahO5cM161tIPtKCCLvxOX7uS2PH
P6sp+WtcPIOnryt8xwt0woXDXEeUV6FRwPzBIMJ9LixSqDEHeOnbyvym6p77pje2WUBgVBI/9gZz
FAtZgaYikxasaQBykmAFQzJenYz9akgCNauOyIE63Iu3lcdKo4QNc3/Qb+vM7hMDD+eV0bdX6j6X
wd5/4waMFvH0mhUVCI4MKvzoI6lhHj6+dSh1QN0UD1d1UYg7wJQ/AoYLAgGSu4nRx6HkdtzFBmA1
2YEl0m5ugUpmFTUc1kD1GuLvl43lKccijC4+yw7MT4vaFcg+Di1DCEG4U0QLNWwbV30V51UwMliP
tN/5fCTcNTGrmy9w/Co6SM1MBjEr7ZjytM54BTt7UL2ks2RAf+iL+lhE8yz7Rvhf+Abwv6C4Tj8v
OVCPQitwYNpUyq8QNhpnjNKGV46SYlk6AYCIrmwWnG25qezBQ/pRUTEZgN3Lz9mEg/aM0520Rtbb
PS46BtTkNLSsEk6JY7HltnHrGuK7ETwPtKlysIvwRkXWPlE+NqTRBRmGNzs/OcC8Qh0IJDEoMXub
I6DE6RTH0Oiri65kRyDksV4JcmX/5DvNP7zPjRZXQOATW/gAnyXYbHDff/u/+X12q2w/3RNDfVzI
inu/s7iJE3J3DVnsTrksK8rcE1MA1Ap6/rrTOgOxwZbfneyHfll6qDG8TEW7AqKL7TjMxvBZNN6P
W/xyMt6ix3tyKEaRdYQipmZo3fdEKRlq/Yb/zOLb7ig/HHzRswpnnlT370yixwkS/8ss3HPlJ5Ol
EJ8Vap5rqRmEaXwCM7LQUqOs+y6vD9c05fuiKqd1+lyS+PGoz97R7b8pRiMfp+PxDCoyLTvcYejs
qyWaf862KTsUIuz2gVDPOqK/5JPi3x4B1jr9PCVI4LDu2oX1CfWaJ0Z7k/c5mdz3p+K/RJPh45Bd
5KyNl0Ub9cyvRmQBspCBD6XpI4xevvjFRBFToNe03YOzRNgBsyghFGy4wgwvGB7pczPp36UH0WY9
G+b84IMI2zTeRtuVYAa9B1hxLhe9cueA3JxN0xLLm/x5QROqHHFt03GXIG3iNNTTpOsxgIbi0kF6
tnsXuTV69Vg1yypkHiaGeBfSD49hMIyBTXKcqtAPt6SXdNl6X5/SSt9nRDiaynYfqP02tFQ1o1/P
Bg2tKsWjT47bvf+B2aJXLRhlL47iocxDSbzWZ4c12tSpSACmV0NVyMwNAFOCFBVdrZ7TICfM3dL0
DBPuHt/+cG6utj9GF6DzgblgVqKFY68KvjJd8GcsjOFpdGWj4B4do4L6qZfU1IteGPPXZr3UOL+n
InC1zHfDTBeu/0MOpmMKGgFibPa4Ni+zmwcB5xS62N0nfJuiTk/KLgF0BZ6s4qU9SYEBQ7ENcWIo
ipjrAv0r/GL5YxjQjmZKx+ced+0b9ANTxLia8W+E79XfQrBmQI+WiOIuCtf48BOvXnOuFIHHTx1g
si9ZvEv//lbgzpZKD0SKbkloavJsCr4L7irUhtQVrwl8NbzyuLHm8ULn6enpV4KlabDld47DpQUM
QplGTd+4n76BJmarIzPQuXdrlJ5YMazX6KodRXTtSIjee+dJ6EG3UAWrmreP3V6P+oWnZmVJqC64
YOFOBkFhV2tQrgLiMalq1IudF7hLbSzViArnkXqlXKFJIZ5xIg8zTppomFl8O0pIXdChqeersY8k
fCDWf6czUMdORKy7n9KiDurQ3wZ0AGe0OlEU0M9amZBwiaaeKOPj6gMUbAXyh35iePVKThvykhR9
p1MRfFd/hnvr+8LiCH+ZwytT9IYLsZig0D6uyvdQ5ue9z3B5F4w1d+PTSQwxXfbXjz25ABWbOp2x
CHlTW/kQVLx5frs4Lq+XGaE0FE6VabQZ3NbWsW+CX3luxlrgk1sqbofBr7hSdZiUVQbyPmBsT282
ub7n4aM9EVJECPXAyGB+ceHmZi2lzBRdThy8KvpkmQ100daE9pfSVujCaPdjJd1hWTEaNxSSlxGc
+V1SZrY/PMr/1URm0YuLEn9OplQj4Q5J7eNj23m1X6kbsaHtE+agie/pSmuemJoaxRd2mIC2w/oT
MWOWG/oSxKBY6UJmLzX3hfwyf1CdRaNEZ0Vd3Dwcak572Kaggemy5ib20Zz5yRbxSxd2absTo6WC
jvvxBeGt+/Gml3WS6RVecLZPMmMQdU/wKXq1Nppdv1beYa4J2gQnJrTmtafaLjDZ0Hccsh1llvw5
BFYgTVoWYIXXtdxoOwlm6lzivCU9PLuwDbocJ2/G7xUxSAoEWOnHc0F+DelVmrc4iGpkgWSIILE6
Lvy7lq7Ml+q5f5rtZPmynxPUK2OxROP7yJ4+SHQ+yGiXd4vWFdCaY7i6+zCgmhf/KBzfLHA7bbdO
Nr178zyxsxdlV6gduZIc0PfjCQ7+edWPCPlclcB8CXBY4V17E9DimXPp1WVrOxxb8Hjou5055OpE
nu7S7xHDu2HgVgLqkIHTfPcbuAhyeg6+eQHXxGia8pJxVveYurKCmlJuX2cMUsOCLBJ+XhCSQjMf
64hZR9DywwYHgRkHsMVbeFUdo7wUg8dHgtWBhBEurlRpfZhfLjSvlkPx2ki0rJRMTsQj2DfTOXPL
uGQv0mB8cgVak60fGsO8EX3OBwdainCiX6uOibNEA6MVmuiRluBatGPjVd2FjDUOqC3Q/nR43X9I
uBT4YJ5dmhxJ7exUepyJm3Zvkthzl/BJAPLa83ip9bcmcfVwou3lTJUs4M2yPCj61ynEN9nZD2V8
NnCqi1r6IznPR7ASdHuk1/fMpE2P83ClVQSm2Z6dcElh70Mt/E1XkyDHqEvBrvMZB+uaSb3kHr6A
vfvraVaE9A02vlWzJZdQdVMBsy5hrlp+10cbNJD15/rC1lreUkuMEOAZHFvymv/ly1YAqHfnm/ee
28dASbKhH8pE5Kv7CibTvCSc1XBCgOTKZYbCs5p37PiS4r4NgF1H6SnBpdWwQW5xdAcUYZ9pClNP
FKl+i329thSH7CTXSrzuT5RZUAdw9R9wBRZLrFrol9ihhyQQv5k1z4CidNE+fAJ6JwlTPxhAFlxH
IVopPPtkMGk9RnIib2zPkkAV3PfgiOH5SBi5zdXjbYqxET41HzK6rjRjN9ziXN46fRGVFw8eBg32
ZOO4wjEABLdaKS4X93xiOzBy4MWgvpMG+33EogSBP8OWMk988Rncv/bCd8ux6u3DHWxni7BAPegk
h9IUkGl/QhZF1qfzD/8EbwNdFrE8TZ/TLj85628O+2fkyaUEO36EcZWVA7vNZlpN+HPEH9uZdfZS
8ZSBy253KOi7fX0vfx1P00o4GGQLf+qxkSTUYljUc2lvE3c9Qgm3WEOGlyuP+HyFkQLIEwhVzLRP
eWPcjBT11TsLfKkEq/7WdF+itIxguDER1wwklpaR9JuRDIxtHOlXzW+XkiMuz5GddG1taoPbzmG3
riVrZFr2WuW5+uaW6jgbXy9DlZUwn7BmCh818OVzqhp+PS42ERLbSmUJGadRgtnnDeTWhXqTj1UG
Vy2SzjX8E0oZj9I6xUprZBefMW/lByShW4RTBQB3mNEOnJ9czWgbPiQY4ZRfg9PhRVdOrrTK93E6
jyjbQ8+cYJWtTUe/sq78GQa6mbGV8xu8PoQNZi9sLloKaiU5iSJfUTvFTI5VEcyDTkFHhfB/5lQo
VKicrZCku6s7ptfVBAkXmetxvWg3REYJ+ADwcuhsGl7S1wG4p3QXc63nnPBYptNcxivJs27BTKNe
OW5KZenFSTUfQ7pxHLz6pWp/JbbeWFeDFzTiyYFN2iIPTCazhG2xMn0KGZicIT+fLvfJDkmNJVvg
5hAB+Ezh+l3pHxBYI9yrVijBdRg0z1bRfWfOyE2UmFYw8/Y574ojcncI2tETFBO1knrhh43unPrQ
P7C8aCR77tY5K7teXr8WSvpqEVFD3mKUaps//2nTNLwfN21kzSR85l6eUW6e883D3lTrtaf46yyE
fazg+6YwGKiSUxr9IklGol6fx5WDZrxw8neDxDuhgGopykjf88szE5u8rEQKfd0cuuiwQOK88Csj
ZyyvzzmKqnEd1erqjtREXxvfMZ3d97dkzA/taD5t1mCHVlczr+JpmydKN1YFk2fXv5fv6sZVhgzh
KN7CU3b2h3zfxO8J3vhX1CoRUlrA4wK4ftEao6fM/w3mFQUHfHUw/D5d1iS+EwMDEGn7C7iuABkM
1WPH1zKg/D3c2cbNwSoShohKYa8Xua9xDnuWLvyY+Yhx0J6kfBhGrr30JgSOJEpkw0gfLSGg2m6V
d7O/D6lRJZRUNghu9Wzs5aFAdZO6T3U675LByxOG4SayGBD2zdvqPqkv8hmetgfRlp1jFV9NUgxz
Zf8JDCVqfFiWqZ3ed2ViuhfBWavUtJc0OjSgQTqaXY3y39rGBRrwX+Y4pXk7BjJu3VVvmVoLYaF3
AQdO1VMN4BXBgFzWHJgTTT72Aj6TAcv1uNPgdZJPtry307ftF8G9s4ECXh0NBySO0l92nGjwjTdc
j0tNEJadeP/v9yMtAUGQ2CxzLx4N8SZOB4dUDI0TzbuK0H1AbR4BHu1VSFkz7p8oK5NPXTryV00T
tbhQmw9yYOvWqb8BxP64xfnf4y9jPFghn2sa6CfLa0orl5cplIWkx8501p/Qo6Nwiyyc5gpjTDy/
IP2SaziC+1jTkHY0R6c3FzuBrWjDXj+6gwWzJl72+znz+SnjPpNXsqZxyMOztT21iBcHN3Dy7iU0
3g5pxYt8JNGMyAq7wHx/alaS/jx1id8mhVcKDPlL+hBCmEXictNAS3+uYHqlZgRtwQnEfO+OZhAk
zAAzNK17G/DFveTYB282MZ8zalKVWs2+7sV+qKBiQx2WEc9L6gtDwFwFuAX3L0CMELhbCEH2ywgV
7PoiRecwfqORMtmGgSzpHJgzpEFY23H1dpJI/n0Ctirnoa6V/ACMLxLkpW5XttuylkCP7d5bm0vq
oElZ4U08MfajcHb6Qh8PZqTS1NZt4LLsEnKZqcITgkqBG0GG+LZjom9neinsNaObLx+2x7CJye8n
Kt/wZKOi2Mr432CrkgayMbAADdCbGfqqJvjgbEC+vRQUupoIPQpeEkKZgh1ctbpZopfgwN3yXnty
nEP+NeWV5Dg7/aUXbk4yTCvVrMgMIfNZg2hhqypP/u6H6GyGSsVXbo1Mg8t+5DGVWd3ZQeBABAjB
ErMSWACr+Ywv0kLMS9EXV6Dfkwp1l+UQpTUjGq68CQjPIjEKds+AluWZ5SMXbm7TRuLkMhGx+shi
znfs45k5kuHbjdfWFUuOZYhhzNvJij7VRqrCKEMRD0cmXhP6/krIr/HyaVWZSUG9M1LO+FY/IhVu
lN8kvD1j+khNtmFAv1M2D29qIqxKfc9Dvm60mN6OEcIjWub7Gydjfm98Acl36Fl3uYnMLa5si/EI
yJJ1dLKWIjQpsON8YbxhHLVJ5seUfPS2vdQaFVUbvKykOY3a3kHrwqZM+789x+g7lI+hIkf6mGMu
gbiis5TaP3ajczsuqRfth3BMjmWRNpc3zIMu4nxpuFvRIlT6rzepL9SubVVR8W5MsZCTCYJVbDyl
2hCvXz2yJ9r/FbvY1IwjpGAm4VKNpMkkGNNkjtaD+K2JjlCe4vR32thO40X8VX/uu52PXkD6yDPr
LgdU6U1HOwZd7xscaikd4aYICTBfP8jiwnt0iZBWKZ0zmED73udyuk6nXAXkFQRrBPUZIIzNpngD
8NyUfN7HDUb16oKzxLhj1ljIBRRDm9He/P2tFyX5YkLsEcUWpCjoNi6XJ9YWzqubUxg8CLWHIAuq
5SXBOaN2+zrW1LQ1WL3NAMifiLUe6EeP8O0rA9BgiRmtXkYyVTcSc3Fo/+tFemMgrZDMW1YoyYYI
k8hEQr3RgVKSPjm56OIYiX+v8qWUB5v40lliiG8Ce3m12V2UPguFYfN8fVQ5pCqYe+e2iXaWgS6j
Ci5W/AzIVsNjiG/5Wd2Yo+Ysn8iqv2B0SUES90wHVlosB5FsLvDGPasFPhO5OQ+2GM9vmi2FR3Ws
9rx9o0YSk6PeOsppUlOlk7Ljg9a4ruApx3A8hZNrStrAKqxexTI32eIHGwibiawBmw3CwBnWgLLF
lhT6DOGh2YsXW0EkXmL74oHik8qxdgS0jG2VZEF0a1E1DDmDhgh3QSJwNtWU1q8QrSLkcGJUywp2
uNQXJqWMXVLB6qlBZsj4UgBYZjw1vrX3YY9ab2JEKqVl8CrMgTV1VgZRjxb53J4eOaN1yQXOvu7M
BKKKqgX2Y2PKSJEFmqBB0gcac8S+B6vZdeHJzSe3ynMFdH9cbE7G2hxcu4pDf09qJlmHK/gxk7vo
J/UMMQIs/rBcIn2bqJ5Gixjo32eYCAbnvLEDs7nPZ6UcjxlsqW6Sli8NGwUBwqkXiKMS2YoZ+Ndq
wsp8dkphIvKMAppjS2Q4Km5sM0dKlVdf1KvXdoeKQphI4zjPtTsdfvwZwunQ1mLCUHig65AdnFgH
HF1feCrIimK3+7K2CeBmk7khjT2zALzYiwlVBpDBKDUk68fz75e4Fghr07eut/pa/GjQ79J+elVz
Ps629PcnNVdACC1Iglp21qCFRNge2qLfsiBcyIw5FNgQfu68f/caR8Je0pPhl9X6POIEKzjOHVYC
26KDK9KdzaZQJcqnBmNPJ5uDIrLO2CEqCXkL4nYqxnyPP+0nAmHKu9U37cpgP93RBuY90eQNEl63
NNGEq+S8HY2RPAAK0RTB/NEWp9K8M8enSQ4saZMmwCL+udtexMQpkQNtX2Q3Mz1S2PdeaS8sCwy2
YOgQaSjPZFAfTyyEdEEQ9RHl8luWwvQnCROTj036QV+6fk/DTCkFs/5P4FAtMF5BdUw6MGndphhN
9hdi5ZonXC9/UsmZfsn+jcH5RPdVYLGO2el0qhn7PqyIiXX0THgqFfG4qacirKI2efRyDEEN0ENG
NI2o6ZOr0yLmMv/92pyD+gaoaAYR5/rYf19fIZfRe9aoP/Aapd/mI4vYD0qPkOzZnYd5fGkIL/eX
HvWdkdtXLUx9a8EkLXVtrSPq4k+UqgmE4PwABQ4BidQalBp4/SDiCef9SlF66xQHpcL/bopOHqY1
fWGasbgv2AjzUdR7rA1pMLFQAS0UYgp4EIBNd7ege2BrCvRE3myjzGkN13CDyaHAn5WNN8qOgmiE
gNnKU/DsJzimwIbLWBUvKD8fh8tRIuFo5+KA1m7Cd6z6KMGGxz8Sa4ZEVro/2495A93aQlyZptoL
+QytOkk+XQDPogTu6KEC6P+CN7ru5Ho7Oo+2n2GFXKQh3qpSJDRxC+Xn2ZcrB1k7M+01bTYMuYLN
g9QRcSBs841pf/vg7yDwA9dBMM9oJQe3WqsPk+SPvkT52gwboq062pQe2C3CS5fbQcKan/ykS4qm
eYzC5o0+Ruh2Hq4BQXHLvpNwv0pD7JJbLdYo+9TprOV+2TozmYU51wHPFnTXVsGMfCb8r06wPvYT
2rab04bvpjnwiuGvmrSPktw68QahmqfOI6NX8uhKN2CHBqdoyVhIRDTS3CZGLNzu0ZgQvAVO6a3x
C6qnNrtMw339S8gpgEu1rik7sfmsh69KRHAiLsIB3yNW8Y85U+hbED/Br1IceoFDbRKPdRsLJf8e
8xuGxL5jIQlX3Ok6MVaaYM2WO1S/3emQsTpXDifjCFlkZUhszb/Hs/6001drEjh6OoILInPfbY8F
G41qN5cj8BOljsYot5X2XF+ume35Pbq8nvIpmpf810hLkgHySXbEdsUkDUTjr1U7N9KCMU/HILUQ
ze8UIPqvv93Y5rXj0vqT71GCQp6MLq66GK9nqnKjsKlq0+uqyB1i6Q6ZhabRS4bbmV5w5aAnWd2L
krdPRtFr3AgvX7ToCD7rMXaBNLZ5ZUaT708Lm2SrYEANsdyaeZSvXRTBtc1r/FM12L7+21e0e4dP
pNFK2suYKLGD884wlWyxvZkMpFTP/TnTiLm21YEAR34MWCTrhsx9jQUguowdMBmLZq29eQPW8asY
BVptzDnuAVf74rIHWKZkSKOLBIdoum1AsE35Ic3aUhxj8AVptSjeO1e5OQMi9pkNpHb3J5RCk7Io
4ZMBYyidqULU3z5MtT4adKR3HSZuHPLV4B0VSfClTfLaqDr0M4e19V7+2rLfx5Qeg6gyCFPicWwC
5OUDlFtPU/71X3cs1BmXC2rQFqljGlK7O+XY6GrsMjzjIDNaTEbNzFMzBmfl4S00OJ1EVOeY8YzG
HeXz6Xeixrp1ULr+sov1jtJC+phMnp0PgQTKG0wRN+DaXivpjHsoqvC1krfbWiJ+iv+T7lwkydEe
PeYEeBHfpNljXNZzaHHbXW6XraDWCGqnxvPi5ApP6EEzf5n5Rd+K06/Rc1dGQCNU9FuHrg9+OMwE
9kA/R3Pe4OXs1fU2yrtoSMep+kvCaKoNyL4kSLxM11y5QyLIbdIYRd0Afa5ktf3ZkQx0qCzbd5Ki
7aPWMICehnQJW/Gl/BLDMK1kk4yu4inb8oafG0y43527tZhgdgoeer8DjMdBHVSaUzJQZ1t0KjAG
JOvEdWjPA5oCFLGBLhzOJYLge7G+plNjDzC6dCkhX+dJyYQLdiqJR3qZuK02md1arYQOmVBJfgRg
V/bvCmOe22hQunerS1wosbjFjHhvvBvzUTTAhaqC8y2kcRhlJUNiYlU0Nyimt2HBpReIC+CqnHVZ
SNePkqyich6sJOvqVLXPYyCsUy/QqMVaQDJ8Jd4tOo1NyBaBbXI/rZv/GHvwhdNcWhE2Z/SN8z8b
O7XCDAUqtq4sHiHUARnfSm21lcjDpHyHz2z34hBqXGrkisNcQNCputYFfzetuQH3XurKAoQjRNXB
hwXKW7dZyreeQtj0icI9lOjGyKwES+hoMpxyDG16P0/uMDiDAOgql6g16rN7teZ1wNdUNfJyg+XL
FOCieplC5IznZtQaECPi+qgAHwHliP6RA2TpDIfN9b7QYKR1brnLHY+yuxl1Jb9mdqzAqiLaX6wD
Oy3XE4nMEDaALL6WGrikmxC1ftzqAsGtda1gGc9i70EyL1EHGnFg1WnzBGjhK2giNuhnihBGhpwm
Ix55pau36PQahvyTinF/nKJ+Md+1QEiuAOQoMlyZF5VG6InNhhiyEh0wVeFIp3lYRu5XO71ej9F9
1IgK57LVLWXlddfw7DvPzYqMQ71RNjem2zYWJiDgAArg8XssjwWM7jqEBbOS6Ac6VsdZ9n6GKVzT
qz4z7avC8FmlBmr/nIhmdc1AZ5PFO8tbKwQrzRjhwDhBl892ll5iQwww6qxI7tz3N0Ig9fbIaABK
WnBSRSfZwL6Yz6Z+0YIniVngdxKGFzCyF5kflYJFpMjEEwbdRTC/I96cXg2KlMuhQ+aNBIbNhwbM
q3vKUsseeE8LZf/N7gydmYJsAgtEvWMi1s/iJETtQAqcbhEWJV3mwZp+yGijlkCH4mmbOyE1TA+F
jd03bxFQOKcuqYTtGbFa//ziB9v8jCnlnEOPBt3rE746/RYBFB4lmpp7Zg9prbgpdk5kjJOHuldg
Gca/s73BWpa2vrV8gLB6m5QpLOjrnw2WrNkqp5mG3Sd9MvhfX2/gAp2OkGbZc+7je4gwgfgA9sjB
JzMXXH7fQZlY7V/5UNDOuCH6dzSA7QKjvOUKjFRfLRRJ9JXJzQ7VHx17KhIRU0YbrzuX5v7A1iwn
rJg77cj4mQ/SOdWBFXv2AqUzR3bHvvzAnHvnpqm5OJEYcuGZJL5MY8iTLI9Lbpv+6VLuuwmPDZqu
Qhu30CaCuFvKCH0StB2CAOXy1puXZryPDuCsrWoxxSrZ6pr4Ofpg6MxkxM342d0TgdPbqvse4/fi
gcwGMJlDkoFnw/Rn/uHTvNs+0cf16IChXE5a227kwLgpV2r8ZL7W5Oc5A5pd5Gs9hEu/3fefnWqj
JJWkq4vDonovXYPmEZKEXWB37c0kjUPDOoFMIIc0/Wr2qgrW+xWuv+7+0gQ9pQZ+tVoNFr0k2LqI
N2tidNBy1+ww2Zz1OQ83ZtI9UlENhzgyR0bycu3Kwkg/UqwuKUg27LpgKZmltYnTHLGSHk82FxDx
P0zIZMRhbkZmnoggh15Nu2dzV4CblLxa71mph+2+lAy6PLNU7Gz+M5C3iM+Xk1kLBUWJM8a9/kUi
xo8SGTfCmSMYRWRVfcpinEVUnFIol4yY420viwvKwN4F5fVaVIysN8BexpgR5mibIj7Lg/E/AEi7
7IBESGlLPQOfPoayyD9xjhRxvMDpDL9cGfEkptjkVGOYk+mx+CPkTOH4xDGIuAFPaCU6k7nHt8t6
4ZJtiBf4/lCNASA1Y4yg2NPlrk2Wni17ta1AqZFhJCeDeJ3KeGd572Cz/H112P22cLj+SkVsREMt
NIQ16AD61VHE1EAhrxBQp4T6ZMP3B3Zi31zfr9yYIoxgTTwVRIfSxLbreG61yLzg54gdMPg4Uv7g
Ozyab+d26JluRKwQDSRolFJigTFX+j2qj2ppfR1oiXjOQ90vMn+sJJN2zauT515L4+iWA5cNaMkY
Uxa1KP9H/rD5LzFBEHWVcEayAAk4ZpZxuBF0lzNXPH6xYdmhSq9lbel+8XN2rQO2s0KZ7gYvsP6M
salm8NZVpHrWsorfL9hLUYFr5He9jzljB/UqZPWDP9pq6rxguOHENR235UPW1D2x5fIHlWTeDLqK
2jzB7Na1rSF+Z5J42LBEbTGTyZVcBI0OcEOZZjUmVKY3s8ekf6YuN3C8T4rA3//QOko7Nt91hz8A
GY9viIbR+phqNR7rScf0Lh/EOXVR4PBnx7JQKQT75UPW9Dga5y8MJzYg928HBGDlL5pGRI74atT6
C+1A8/S5mMZvTymIX8XqTZvCyZ54w1VJXkyP5LhNlR682BzY9jraKYI0kbXy87v9AGGnVxvD1Gh2
LOI/1HAw8iqBl9UJQaxdfLSK8ET96KiYb6VXuY0n8LM49EXCceDL9mGn8TXKQoTCImWswUgJPT8F
ofr4TrvayDOrZwest7Z3gJFWrQCJtCAMLr4/mobwQEaFyRoVwZxSb1CvI5SQz6dZahvDi4CRy58u
qrg6l026Cb9Kz8CpAWs9zzO2BEDqYUlyhdjPGjzG4MdPpQ7nrR7uWmeE4jqlutZlc8V7O4iffVpb
VpYpb7PuCiR3gsj8pnmIyLcNUWPEnFkHq69yPZXe5ZXdDq8rGfMkOmvNnC3h1HWXqUTjOYq+dA0d
TjQi1VWDMIH/vIbsjpwWtG2SqMoUKhPXhu0To84O9BYQQppaRIO9bcfu69J5iGAO5VI8/8XrG2uF
u/HHvfPsFuyIB8oIV1wyBloJuqSxESxOYMgFmsjpkNJNpVABBDBedogAsdFgeZrixcBKK9andtd5
WPxW8HBvsoO+19TpGT+pHRANarJiiCSwzmK1cbsNvmw2AsOIE9olwmK+y4eesH4B5E9Rmeys4PKp
or7jra6iG7Lwatc/Y6H6wLh0Ttx+gbFU53pP/PzoX+X3lg/XK8B3M9L4G4UHHzma47wOn5GQq1hL
pKSbzCjIhP+1O1hygiKZUJgMxr/AOxwsGrgoQ4yXbSielS50rjZIE9T8S5u4xyw8wXT+SpPwO3r1
L0OG+ABK+WiMU+M35TI9Sl2pMUqhZ9hra8wivlLHgVlReIuRy0/s5EvOtspmo9t0FPXlsKlHrfZ8
ETtMyV6HCmhyeNGb9PF3xb/ErABQpawXZmQ62oq79h83xYyN6r2ddUXTwK2oKxCKSaLNNh1L6fvw
j36IehMTpNuCxHLaGIm2dctU6LVsjJ/tQuIvJFzQBgv1nB54ZLwnDQRH8xMp8XnKjlOfE5OsrJyQ
RfohVyedcmQpCDQamGcsPDFE04Y5DtqCTTW6G/qkYjmyKRfmzyfEUNmSttD2u2lsxisLGfGnf20V
52LEZ/I3LNWh9DPEjJcLQFgl9LuVumLxIP7oVTjqZ9pAlTcrtPMfaUNjpYqDHt2PtWneik+vUKka
VbLjskM/WFFvJOWlYY4MFFwZQB7it4sTI7hRnKjmuAgvQGA0PmxIhjCt+EHc3+rxJtUvi/3hWplq
0zmURG5iw9Yj/qlyBpMqbLHmUsqv1IV/kjvKhthZBebLIyH1GzdzGa/iEPTnJQtRMZxXHJUuMEtR
aqa82ZYqO19hnfSCGY9Xr4mUMtxNZFxvITs0B6z79J/P7MdslaaEWWUXc3cCXABlD9wqMh31k0Q7
vSWI7f4l2621gdvJ/MJqZ2KKH0yLan6UR7/A75BaWIOamUbJ/me0FLz31TraKks7LHyS+RbfXAs7
pzNw34fJKk9E5FZA7xSNnL3OdEUlNFPFapQEIK1EvQxM8mTE05x9v0sCzQZWLXxC6xXLWaTeAvY1
gQRT8598ARAbNRvLbTih10H3XcK7E5QEmKgn+K8pQy3TYnLU5+srqWkzOUpoUzr5vg9HRhIf6BO0
aDt7Xqpg38fXc+fdpQ9U3G6ifVxTZs7fXwkfmWaHe/0LaAGpFYzBw1Kx4Gbz9KPQs+k6fk7C4pS4
JS25b35NPlUJAIwGFvPowNNgnx3mZF380OhrwBg1eT/NY03EeTrNNTjD9D5wDADLLEMolM4PiZxe
XVtXXgGI33+edaL6mkREJa4dvu1meWZ/0Rg/SUFkwheD4+cxz0OnUUf24jMNFQ0qpyXYC+lazHDs
MWhSy6Wy4/rFLKa6eKTnmhvJjL8YF8SP0gLR3yuryllteevW77HIQHDAiSNbpCxuyjVXkDCyDX4P
6YjbNbHwHcUAwo8dIjS/RNvdFaYrIk1vVfCyBOHqd8QOtcdfDJhHjuzt8INhIL6a5kSRouL8nR/W
p+yAGygTMuCuBPXS3p15OhVxjnZzidfoQ4YQGwL+nm3LIOop9LRPC6PMSza9qEPNSvH8XT+009M7
oVDas28SllwX/17eU2YSliUzPV/zfa1Avz3jPUXFJyWpwNtk4rg3wY9XGCa3ylMY7yyBmrGo30/s
Z51o6Jg6F+rG9KXj+x0JSnK2zHISfWk5Tb+uF1BzQBv7FCGdLx/BxgRTIsTPE0GehKDWU/8w3Gkg
SHArFB5Z5ZRrNn5qlz84688nDQKiSZ1/DvXSBASm1GlQQcml4p7qk71Uvu7/0cGfKDxsRrKxDMrf
xxZ4WbIw39yPoAngyFx9s+xSNa26EAmxf1ozjvPnoIMb/zl3iJzgHIwCiyH9rZDN9zEQ2JTZSPgl
HR6ajhasswlS/zRvMIh1XIeTYpiLqHz7EOzdBpdCe6zE/1UpAdkrR+Dl4qpMQQYsigr4h4CwS9Qx
A1Yqa1rphhK8iNmgnnQX6EdBAt4w8gzqgMJcfQnmdsVjsM0JmxG/Cd1T5fcjh3Oaho4JJxVRjCQo
lj9/JpDVobc=
`protect end_protected
