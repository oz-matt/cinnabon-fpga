-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
sbSGmTARFwKH5p9nidlZv+qYTUDLlgf6K/QY+GAK4Ofwjh8fYsuW2JDBiv71xLhjdETFIHkhfNDx
J1T/SDDt1p8f6kgDyK3PmmjU1x6XLrgJqogCVCjEGEd2GZt0fpWsolGiLquS/pCkk5ExCW86Xoe2
0iP0PZes+3rWzs5ocqJxsLA8vxLqIaWHUEQpE3idQwyzAzvmd13cUqOm/F0ZjMzz05Vd1TC/+8+l
3VUJ9edi5CuAJTBYeCeCl4E3AeRDAX847Ug5k/Y8E9WSRTzauJh4JursRZA1h48LzgIQmeQ3jdcC
b6HxdL9v2zrnDgdDGA6N0xVd1E9lwpNBKXrbjw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23968)
`protect data_block
qLlohHGQW1dhaAnNo2Ix6+sd5tcpSVLhorH9niTSG3NyiZvZxNQYo78ss6vNXgNM9uIVu2jgZgQk
UfMeVWevKgDS/JA0oIQkHcHiiKblcFfu467ZypCMRZGPd/INHJqnMUhoSVlBqZ+LI09sipMRSdal
HXPy5GeRNkAdOUWMtvQJlTt5/7a8+lv/N/ffQW1n0kmT4bD3tY2JpyFkdTI394FihW+dqmExeMX6
wUWHjBfHXxwT7O3CRDjps7sJyzMAuHMxIlS0FF6txRt/ANxbSFlmm27dVr3MqgowNPhoFvj+RKs1
w2riVy1ONY7AE2iLwBv+NtFm7wUWrjwwy7dPCXnr1LKcxk+2V5g9xYJzUOwJZXHgAQ4wgciFcm1m
SoKTQo8Gt/R1ultocRilJ9hNi+sPOru1F05iR35zxyOhMCn5jJxKWOma5UziaXi0vTVkmTcdUTFm
qU70BL5heMw83vcH8Qkx78/n0Sy9VbpfaOJ5jzJv9sSMsD8fDn4l8+L9pf2yXTv0bqudylIkC2P5
DHMI45tX9NbgCsxy4neOnZw8ExqGaBxirHM/Et5cvNUcgi7vFUi6iT3aY6FXhS+MkXFgA/g0uloO
EvbNlMmsGHQhs5k+OQYf69jQPfMXn3qiC8ne5pTnmwKFVDXoxy4NrVtzrBPTqdeg/GTR+GQJ9BTC
ZD12UQ633ap2xeFGwaQzUB9e9VYjnvIV6TREBlh5AxVPF6PcfqnDBDXCzAzpWxSwn1xrlClihV78
0Qy8LJCcXJSd2YgmAhXK0kGhASpLjUA5xRLxzCa1dPXimnCaKYmgjRDxGE2M3zdVI6N4C2a0IXtj
9/LDPNTaGjlEBe9Tw6gwglj4ncO9ISnSZQJI5Y893htyRcc0ijDLK44v7E6xDDj5MUZyVvqMNOkw
A2bkRWFqxdU2cqibEtsWWUdpJWRafZlHXmDi+6TMBwLT7KnORcSqDENIejA/1V2EG1oBOeHeVjsV
eX8w611wyusFiX8O1dxSiljgghDyD1820JlU9W7L5LmFTEmXa58OExg3ToDbMvJuiat/gRN/PMAP
F3OFPDOfA08JBdkEbBoessYVrJDFW4yatPTDl0qJHsTCihHSPW/lE1gPX0mtJgBJFAL8xq59tzGB
uLqsJ5ofmAFlJLXygQGb8PdRr/8tyiCxstaoEnURzcks+my5P/t9W+a+FMzRsZvS+O56rxleF9GK
0ysjSdPP72/Doz89iDJJTcaUirRyvxSflTp6uO2JBlyLj0TTuFAvVTs3Q7RX6OkexfGtleDhnYu7
y+GLMFnY1C9OO7DyxJXl08XxO71l9Y7Z9XOQ7FhkKY7e47QECUtzmCfHkDGBFzuW+Lt+r484zVLD
K13dy+dxVto0p3n0eZqiiWOn0bOiAIFAtYLKhrNSL0FRc771tg9GW0u9UQH8pYRJm8iW07nN6jXq
9+H5Zc4Inb7UzSkbEwpoxmaqA6mwSQVB2FS4NcZwjQw6Gk0TafDE8t+6QPsFasj+XTO7y80RqsO3
txrzc+ZcJS1JTGoCqiHjqeVsAyiQAuDbsNVm7p8ZGc3CPd+TAp2c26Ma1B5wnOFNuAmvbQ2XgYt2
pBExEPRAknTWydbtgkpCq1dwMdVnK5fLBxt4v+c0htYA0qNciXyoR3wPgLxl8Fc7F+FFuw8pEyOr
EFnlS/3x5AZEeiZZ+wK0xjRwdunK5frwQKMj5XWTTEBohu2aD+NnYiLpN6/1hQfn8+4oUgbPK964
WpEYfEAp2E3bJglM1GFFhlas/p4AApA0TRFT6b2M5VLAK3pbOOgnHPwlNpCHESG5fNbeItphkQw6
rppjN1ZEWKqliLDWNu7vmLOITwLAF4VfScZcxFTLG1LOkMnmiK1rLW2d5q2SQ3KrywQWiHnVqoHQ
l/uiZlLqzJnaONa/YS3GyEWJewSKt6BfcPTGLsA7z8ikWVMN4MMgqAIwT49bGJQHfYsbMKhIUe9a
SiSbhK4OyXpGGctpcu+I7affjz0CqirYPsCPmuzHNUNPgOH6jl87FwHY8SmI5MPRWN0s+iiD8g0Y
p1/rbU4erMNHnJhhUJzrwvFLT9p2LeQK0kO+DmbrNUBBySY3LsbBPQp/CuyJ4y8Y7bAZabUn6j1B
AkE8uG4yzxsVomr8UIdaTmJvJVldqFbMpQr/hhkn+57G6/eQTUy9wMd6sRYG9teuHCOJTL+5Tz/V
6gFqeVraY7XZw78lJGT2ESwgw/vVB21KsouUImIojYsMNxhdAns1CSHOIHjz+ljBGHectg6DO1Yk
veyMvnIBtSROqTsa7bVba/iRQkY5zH6BY0yUp+tIxdR5YXbqHewgsgR4qSDYZWSQl/jQjcsMU5FR
MrrXDonjsjbFXLWmyVKiv1RCLMUHCdrKFy4hX36j+wwL7SUMysgh/fbo/iWyY1IQUEegE4h9aybY
PNQ6m1m/uGpv/MvLq+SxmgB1j9D3XCqDj7dKUT3HEQ6dEQI3IZL26+14UugDTnMTVnnS7Xz3iBJw
JlO/94FQxftAumBZQL4YuWhiu+ibC7Hpcmf78p3wEzk9KyKhWMWiwh8I6waNior80j4v9+xvyY3X
yZprHLygtwMDR2P2Zm1jqS8KDzMBjbzM3JeCJbVymCglrcZVD1XJRy7dHMaqBidBpF1CCi1Abvhj
yEezkk4JcD1BzHcE2XgNjBy/iZFlNCQwvfP7WfH8v9hoWjL4xZ5QTfo9ki0TSTY/+TO9HZd0+b3c
4BTuVzB5EOQzmKp4mCBxaS0azS0XxO7ODo64+0K6EVyDRq6P/jaQU6gKjr/778GBy5Y11gcRBe2w
V8snnph0X74ZZMDpeU3P9TA6UVf3djnCxb1Vc4VVykm/5sWrMBUEoMuvqngyJWN3l12TgLUM7zhb
mfkPjsxL1YKpsqdOPHYL23gUPzbmepjgt8hzYpJVp+kyxsjGDp+r/aR+RPlZEigyTU4unoWN+q7h
1FvBPONwJUTnQxtAa1DVPS82TYJLy0SqankjwY0U/vyy2K8We6acgfm4eV2T38ycK13lhKHp7Yvy
PrHCAiBkYVeOxqlTDHcsHGNXrJRPTEOa2bQnzpss4S50RcfW8LQn505egyR+3j5xD5D+KyJwP67n
Ppy3ubGHbMWutmoYmodxVSlEUy3YDS8Mw3LPknznebAyTXY4Mh4tT2y7jzpktVlfAy2J6HQDgLgE
71V+5jSEqOcrRe3CO/0ReyfXpedNax3++yUDdy91ogyYKUXLim47nCwwKm/Kqn2qx/wnr87Ma22Y
wMKMooalrBDi3j3S0vrjvwS1JhshfX7+kl/kbcIHBeb4QgiY+gGRf0zQGCQ0wBehHJd5bL5flU8+
CUZkyrjTA8AWxmsQBXrki3p5IggcHi1h/Ntk6ArhmMOOggiNSyXyE9eFLBR+tRqNkHIIuOfWAVAZ
XB7TUBf/FeWN132Hoh9MtuFIuLHXBbc4z6wap1DjwnwU7r2vhdWHNrqaq0iXqSxNWt8l263ztP1l
rnVmB0qLbYTTkYbn7p8uYg5Ud6iYpPbLrCxtbHkCmDuoRJX+F0OTU2hGU1zBrt/oGx5tKEB1LTde
XCwjWrj7e8AE7y7KPwGn17mHz5aZu+oPuPfLuvr51S97e/xb8pmPVjbgm5qVZEiUw/gUchPAZPX7
sKInQMHLLe+BPp9Svpk4LBJQxw2ekTGcQIdwPZyAAWWV9abt3BV4uFuT8nXGFDvqB+UqJ+uuBxDH
brU4R85Sgyt7Uti+u3/ZV/dNXJoUNUK+Faa6bR+JVGcabJkEReGW+OK02g7nftHfxjlmTk3cz1EA
fSzTqcK4qO3DUePLuI02o+sb9PKVw8WoAr0J+r2tIjhE0v+UG6aU2WORrQxXLqOSTuxXTMSs2lAF
5vGyTIAgSZmgMHShtShXPrH9WegCtw3cNb2V3gzUxpnjg25+3LVCQ4KROR9X0EpD7523jUjNUzwD
N1muJTjosYlOF/3nnSGA6sPn+D+wbOj6fyaJokZ/djaSXUDHeE5eAYfzGOOjmJ6FlvvThYRIieFA
Fd8vcd/vt+rwdb+l7XGCC3LS9/wcYdLAzoGsKyBnsi1I9IEpzVzqiDQDFZ2Iq/hQ4PteidQWmiRL
40F9ai031cZRywfAsncHCqNt7Z/6OBA/BpQ+4VQirPikycwiNwwfol4f2wNb21VBB1hbe3iXSZyV
npRvocw5WnZZcRNtRtVWCXz22AKRWurFNhHT6XX+Do7GMlC75dK7Bw/9WN9YBHxZT1KgWf4IBsmU
dcFeWeOAl1NGj+cA4Ruc70/05zT8PQwZEmAhVsAmjmu133+pBXYxOpn3cvTWhwRaQeeAv8DvNy52
+lD+ZhC8KtdgkHQPNXoAcih7pxCJVIrylOSilNJ1r+0uTRwfcE7IfFKW4KzLyJW/SksRYaZRe5FT
7YAvW5WCuQuBsJFNrvTAndYPHByVfxYf56tCRKVMI1+IAJVA3VSGVij6/KrjBYHfp5p/obcwTIJP
neADqUKr74bEChUuge6k8t7+Wp6vRhwkimfaDI9/pq7K5/+G0Jg0B5aYbAXeigcjjz4sBOcniw47
nzyqGA538oPWGZDxdJoofeoWLgzL4DgzhRcIdlht6bzerXnoipD8HoVDQqoyMkqKEJCon5z/yRzE
Rmp/qwxDOIiHaBEW32Ekfum9pgksnvuW/RlxVQiZLVwkWOhTSYuiBiFaNQKBCKNXlPEbZzUUOmSM
9XsuEjJ025FTwMoBcOO82yRBJgzuOs85XQCvouhOCSsxZZi75ZndW+eH5CJeGPG3kVyhSAIB0OMc
RYWZccxFlipBLb9UfpRq36IHCfW96S+9TofcPhCWllKNI4+huzioO/fHoRrGIe44aA6a7Op6sntQ
YoheQpvJYcRuFXW5j7PMbgIthi7rc15SHIq/1JUDFYolYQVIjw0KFFWVtU2WjvunoS6HS6/UPE+c
G5vLSmJ6Qk2h6Au2kpLe2ztwgXlClpTTylu+BuUNfWHiQqQxEzKCsP1nERdP/vuqsDeQ9uTd6gSQ
mOjnOI+BDf2Mj1iZgYVCgwgX5s5P3YmYtTwCiRqheLoQqX3saWG3pFhPn2R0W25757dgMGF6qvTP
ovCjBB5qVeLIUfIXuw7Gb8NZ+4JZL9x1HjVXRtt8cMtB1045+xxfHPwGaaN/amL5Zg8EcOwhnehL
i5OCgniMGMoyDwBmB2EjqzsuF+bzFy3jJDCutv31kNRsUkgUb6KoHSemXqYCdq9VF3hPU67FFJMz
/mIL8Pa+6NbJ+FDAheDjcSQDn9Kp4zExvSINu/C886HW7i/5Lhoy1qTxaVtRoV5k5y5q5y7Wxg22
IHq33jyoEocKLXVYhBCFJ1JRNDO9c6zFsRLidCwlaSAi27O/ZkiAjbAOx1QlWdabokkwqamVg08A
RBqy+/gStFLatEiVo7nBQKvroJ6M9PJMCQkNaVw8Mou231nHmzU0JGwNNIA5uOG0lyO3wyMzVAsL
oPYYgTi+xAIGKqDbBR3MEf4Yb+4yOJLg1yJgwoiMzNeoB6/tFnl6czDu2tJsNPNSBdkLnwGQ0OOm
hhac578lqbK4d3qImFg03hhBSx2501whN9gjKn/FwldmGhIuhSuTCP24J1TsExf1kxi2h1+/VTcM
tr+CjqXCHP2TNn5vSXeOZYfwR1FEog/lJtvfHHpCuk7m4tuTHUkrUO5aRHqEqfoYtDbg8UB7pauK
MMWbEzys6HvR1RwZNAMneiJxwT2r0zXPKJ3hC1UUFctnnErLPAM9G8aDqDYWwjDC+9IUxVZoYjmq
zKb7sni8GFez8Z8dc1yMKcTNrzoRoeXzqsXYVlA/nmTDjxo0vjl1oe7ABjWILjTnrXjVu0i6w7xz
Ps3NY3OKZlUfARfIZMiDH91/yP+9uplZ0Y5GkMFtDHtRJ8jDGximXC4ZKB4HUl+Mv3WgJj2BgQdF
tNgHRKI1YzYATVvbQg9pf/yss1igyvf+Vh2Lu+jKqO99l7iuEM1Weyvdc80arVnE5tgmm7J67gqH
NClH1rb24Q3bgsqGb7afJ5q7iil3MegPc2zfXmvWEf7Ler9/+U7QOy0Vr3xbFudgvUnjD+LNKnDG
Fswj8vy7SUe8oghVdS3bodjaKbauZsi0keBlsGwGwubdRNUXoQCqmOYAZQNgoIb5EaTMh0MYFFFZ
e/izgIg/+HEGZLNk8LX6k32KK5WxtLzZCFDQiqUrfp6L8zRgNvgk2zljDXCxCr4XxNDNIKA1USlE
bqRxqv4YLcz2Bf4u/fXOWoQRpuQUYLzQLgiPoBYAXtCNELsbTw4abQRZFE5ggd1uxR0uV2irFv89
Wj6wtzzoXcVxeLZNQRVH0yCJEpVHcW9TW5reo1ECbBM4SNq+mVgUH8Dpp/0mAgsmpClqlNhvAMMv
hXh8lrDsACm24w1/r7U4ObGBoDqcU2/UW0OXmsgC5LWBfIfwOoclbkHillytpShknsOiTt+WZeKF
L9hjD+MMtIskF5LFM25a/ddd0575g2Kwn8wafqpWPWtmPkVozm0UtGF5uem7/xZ3yh56k400txz1
IPTrhzlGV+Jwji8+jwgWBl4TGVbadU1IKbFawuSUzv9FevVpcPlcOQ7RtSxO5mNyF4rhRNBcTjhw
afCHA6NcW30mMGy7tVOVsOMXVXXu1OUNZwaOWoOIYn5/C95NDlIphxTc3q1UjsObm4TeMnhAD0RW
UGMgltEnnngS+m362GxvgfZn1lEzhpbcOhFN9BtceQnozRbgLHVoZ+8qyck1aHn5Ll4ZWsmlxVNp
4dMxHhU7EBD37jiRLRhVmvJIyfDIzytuNAkoo4ngHCTgHIjfG4XjjM10B70hAEPrizE2gphazw04
irl5f3cnovA8mK95md8WHu2DmIZLUcWYKhG1GAJYEH4scahFNEFWQamZrEuhHt/WPyFwo9pEXO6A
f8lvhEoUgpUr1kXc4u6QZf7yRrH86dwhtHEKobsJuPR78RGfN91QvJJixMfW0UZ3A8fpvUPAgmUv
XnndxdpDjkJ1A7gGViAvOtiYrnDvzr66AvJA5tlTA4jQZI9l+crPq/gAXaFk+xTAIrD0iYEra71m
MdzNU2uU+uN5PAj+TVgZbA5TR/4uzkEvaK7E1K1aAlT/tCs9+VSu5UFunZAPnXqWpTOFacLCm72X
dLlcavKPtXRLH0cnBpGrJrgs2tqJIfmP2onr+P0iEDBi78DQJ6P0/vU2mBHcLBoDP9dlb3+YQDGG
QNFdSmWlRzmweRK9QKNgBFalucbtGUwSU5UKU8JLZhU8GmQq1phdGdkiBSX+BHet8sJe8WvvcaKL
xASx+naVG70hXtFArpZgQzgdIubFI8AATWJBUgmflqs6e0djCx2V2y1CcRBPMAzx8RkMf1XoadNJ
IwzBC8scyq2hnyiYJoDm8eHlTd9I9ee7j+9F+3JdiX+1uSblVHZcC4wojGIFtVads6IUSGsvWvzt
wPr3Q0d9oIGuz8y3mczNI9IO6YHBEJtObjwKa7GQvBRn+MA2LpigQ+bTp2vtYTKXRjOWpv6u/Rd6
6gc9RU3tDz1JziqXyjMOTiu0CsGTCNrpjKgzcovTO4E+nw6DV7HFgjkV4CsmDBB8+KzHwNt6cfVP
9UygfJnkAz4oFGziu0bcxsKJY7NkKEIH9TXsPPPf/8cHZMkDxz3jbd7BZ3ScFGroOGeKEjbC7vTt
noQkqpEfjLaaP18RAIZsomzX65oJEGgezGNx66D7marf7tPaVdZAU1+MvI1Lj+DM67uwX26PHD5a
j05DcNsaz2Xul5An5Dahy7jwhMDkXECJfVIhpWhEZCoy3c1xZDUpRcguUyeP/fY+PWSuDNUNt8ey
8kcVfDyslCcoFZAPD1WoA9JOaL0FNjxvHoqE4bSbIvO0ojPhAKtxK7twuaTdBI+o0hbwCfY5pjr/
quGazPNI6Y2fydV6G9XNWOQAXOslMmRxMB+0hbzU5qVr4KJdGI/10PdljjW25ep8y/j9qdOfxAM6
IGi/NAoj7C3yZ2NdrqqQLU9eMWtjyNZnybp5IFCQmzVa94yZyJBXai6fpXrUU1NcBpXUvRCriw2k
jmPLutiqw2b6ldhec/wBPZPCQEUzOlQml5lvi5WwzB2xPfnbhQcH+Q8znE/Qj8UsrVSTpQpfJ/in
YTjKTK8THVvmaby0x40MkY8iOMam1ZZf8nscMnG2uoV/UJPRsxwZl+CeJMKH0+a8PIS9a+7IuPyf
i6b23y8A8nOOIMEyx3CP4uZ54JlH1Bzg6OM+yxDu5NNvyZxRbWBbLr1eKGVXSddWmRTXCYT1wwSh
kpRo4+PMPzGbnz5YRUOOwT9Xp9lz07rJE+QN5Q6LkU+NPd1+ZDE9s2HwPuvHZ6GJbkl6VVKy/669
/KU2eqoyhOUCDy5lpgHNIoo6oanKcAp04zh6ISeCKVpuVTjQN+N5Z5fhszX804pdxguUDYs7PqQk
eCgacaZ0qakj/12dAp/eW2kMUa/Js7XfV0SxHjTdh+prWDHXnNPRbt9fY92LMU2AUR6zEQ36pLxY
4YaByKQo1M47rZBmw5fDSEQKgfhcckpYSQEYUARtwwjJyQcVtk2uaeLguGdvZCDrqqey1qN+TciF
RlS539xjmoBUTeeBz7jVZMeu+IbyYSCwSe1N/vLzHD2oazp9j//4fXQYAIcoUe4W3xnwTccPMaNk
QDXH9vGa/tax9X0ezk4H3QM/XIdGL3hERGSv/mYcrwN9EQnQmlEc59QrZnKKeEmo7I21ZDYPSq+P
kh/A8Ww+FSmbTax0Qi1GPdgIkX7ZyhQIXWMKcLBg/99jGKuUSX/OgvkO1J00CDu/gBAyzgYO3ojn
MoJb1aae14r8s9oLNzxlIBvCOVjoYLWZPoCSWkDJ89M+9Pkc/QEnA9G6SfAFR8mulFR/AbhiH87z
OYHp8ddscVq9isDmcpI6hcito+36YcRTlUigNHqIlg2lGDHocmnUNhTWwMP3ANVmq+rOnRu+4rJ9
V8Z4aDnj/XsPDp62UapzL0OG/hZd+VrzTx2gzecpp8gm+QmXs31YjuG7Jmn9AgHdD3+FdGyRRLQi
9bFeBb5vxxs6J3uEp56hGX43JA2SDsdKNNDis686/jHp+m5B2M+9px1qpOBKJisto0buuWnmBaXa
6KBTvZcsgqwreoQgQB1+jqI/Dk8iIAnl05sRqIlr7Uu1psEKFb8ouyiJ5Y6ZgX37go0/qH911xIJ
BQqCD4DTCKqtA7HiAE4vqSAO8X9L6OS92RGanzf5KOlu5X/L+jWLOJv5dZVauYDKRIpO9gRRXYP0
9f/DjK0cI0d8GdiKPTA2kle+a6oDaTgfZ1LPwQW3Lp9rC1aBLW5U0jlk3l/yPJ4pzKJPvfv2jTyx
uh+h7jAJ+Va267qB4iTeZigz6/eHTadSfoWIBYVqJjNYzL+IcUi47TYHlIBUvzA3rZSxZiRD5bEx
Kc5KpVc4DeesVyhKFP2ZuTAEEsW3VHE1ONKnJqqR9YOM66OkUpfopr3fuq3q9WcSjk6+TohmWjaP
Yh/g0TNClTjqYWwjTsVy4zFjX5vD10SO1RVfgwwqxvjaZa8uOUggCvdWzNTAuCx0Ft0W/Cu+5TgN
Ce8ndhqkio6kV8uWHObsb7+c09FLVbgjXDMG3zMQbNQ2NEcP9AK2/i5kPJ8iZs21xKUsT5pAMGTD
kd/YpuLsf2BLOBPJ8vSBZeWEcfOX3BRE0mhZZZwiIzx4IXSRUklDF1TnSYv5YzEWQ3tGjVfcHx9A
qvdppN8C/Cbg81uvOAEp4PD5wxWxQZygKLCRXR6yZm/MhbeGTUGuo8nf/d0y+07tFLHSair++We6
AGPdRt0bMajSIRs0TDEKxEgehziTYIfMOfhwFd2AJQiscDfLnu3IxeVjYTh3q3eHlUSwKFuGaRVy
Kv0gj75W20U68zjx85GtEH5MiCSayDnaFFbNaJfQj+HQkBQOyPD+RfCe0qYPB3tLZXkeknGLGavQ
9nyBKDGILdTvJzAWTk5kKwtuX3XbTSj9eCxHDRM54iZvhFV+DNDQBaFPQjYV70Mvy0ocqZxgjnNO
fVZ6FwaSuT8zDrIH/6CCCCfLOA5WHNM+FWIBDczNmE31TFV1vBi6uvcJYjz8D9JmiO5RS500IEcQ
sCZ2A7vfNdGmaiI5/LK+EQ58QFGzmmk3gwz6EDLca8vFXkzgVK1tKhpi5Cdhslrl5q8Q655u4cjJ
TFnEaby+vXuwPqYnw209hoN+Z5xYR131inpndaUKEy3xYqzwtxystO6fpAJ9fnkk/Ahiy/KgS8fD
TqioW2LR9DVqpaMoniJS7EQslK2E1rT90sLLsa0J5wuKHykvv7GumXRvfxR/2knUA6TTwwcXec+N
aePG9HZZECzQ+th4aVEXke1YCQrz+Ix6ryE23HtHT6ZHLKZ7NjY17OFtf7o+Gv7+Zs9JLGNE4Z5e
BIVoQbKJ0EbKdF75ztIBppyu9KzE49OwdoNfviGUxMHzoE4L1pukroGnWSv0BmiIkSy/s7/OeZpw
RqQjckTo3S9P5z4ziOYsUUToqW9H64WQx+RTDx3ZuDPUaIKnmM4SguzJtT79p9d2CKyFLN72m11I
36WyAIANP7a5WdY7TJKpwqt6Slb/kXp8MCuH/OXnQmP03f/Yr1IqH8UG5knZbfvuHPy7IWRjh3wG
xSm04fvY5Kb0VyezDaV/bQA98v0kApsdeQrwRyFTWRxhWfDHeYnBhg8XmdefOnOFvFIb4JOakEVR
UgMXO9OELFCshoZuZGyoZtonO3qs/ZA5yMzF7QlQic5vwcV6DqWD2afV1rg6t9dv1vmiBwUqBdfG
Zo3NXwRYkaiaUgDp5cXoDgOxm4RlvK3nCG02FF7/U4VWgWEEcQfTG2/hVs1hTCPkjVfQG0ixE7aD
SRB6eabLEf819bOpxNgh6eS0wdAZdye5kkm1sfHfHZ4xkEqT1HsE4BAb/kN9Npt2yQjgkm8xMKZB
Ueg1464kB5FIJXc2CjcI67jkYgrQD2EPv6SXNxSTZcRyWII0dJne0PGcX2D3z1HsrdZ+z/g/YkQm
W8BOXH1oQ7L0pewauulJ2mkcJ5tpATrr6aMrnoKPqqivG/n5ebeFRpiFg5T+P+lCIyvt+PP3SHVz
ZYn+tUVvMRS52d/6Hn/PE2oDTwjoxDZnW8TNnkIZ/uz+3ro5R52gEvFXNJUay2UurBt0cq0X0sbh
cQ0eqkHdpmXU7pTulv66cxITqIkXON0nG88fYMwuR8wpyHaMiZbk2YYRzUM5zIkIFAXO4Ob8h3G7
Q1BmD7EMeM+EJrPN2vE5ZbLi09UGnoa4YL1pzSWNLdyBYiklZrXgWLsqMBI7T2OnOJuDdOoGp+2U
Eud8233oAQUVyvb3sf7X3hXHWVlvSS0CQ+1iEBoqEW6YUBMdC1x318e4QCKoIczS/IWRfKv+fXfY
BQOsrRTqSP+y2ryJso/ggMXg97NXUMZXWhorQxfOXz2upNArbwl9mQCfGDLQ8GI99r4sryOoqUbE
rqh5zVVMad8s1Xtf0mjYOuPWhov5LCRJqJGr6ns2Nb2RqckWc6gBD+tIeVr78TjfAWXB924foFpF
xm7YlxJNIYaq5puFLa3d+33aOuH7tj1GhVO9H5ifUsPPc6kklDpBo8BpCiwWj+xXC6U/CMeRyKPn
wfevGx3LmQ2UmbdSSK1/hMGh6s49qq3T8n9Z3YlP23PBnOakGyodq3NahHjjVdFQCilMQ2hsL8Ub
PhS3oCkbnuTY/euI9lSMbvAJnNIv5G2hJ0er0GAaihTQjtGhv5YCBzOtuTJq7k0c2AZPP8hWSmtW
aDld5zqGKxXR2AYjhVRpm/AmoKvGTaTJfw6UxeJGS4IoTvv0uvvQJs5gDi0LzRoKB+tImimOfiH/
PxVc09aZzboHXUOp2PRmhZX72/DaXaMlvXHDlQvOZKimn2oH1z7FLiXdI3b+rtOKKZ6m9nBQW7kr
eY515VdrxtESpn4iQz7djbXgWj4aMvizZ8BoTCOdFdvBu6sAqMsIR9hkOt9QHWds2lEKLrN33uAY
hoe432XcDeljljYqwF1ec5bjBGFtrRNEtHqzgoBggEYfvkziY6gWntZ4nedIQJVjB9ikmg19OoMB
YcxaCFybFrQk5mfYaFnt6EvArudLfS9p/2/Zp/u966xZ+rvgyy811svh+C8+mBliC8dx+nnayAGT
coyyCMXR1wUe60ip7uOHUzZb4baM/RLG3BrvC5dgDuBCsu12F+sXfK3MGzucoKY7/PHSEcmHf6zm
YtOBW7PdV5BVvV7OfHN3Egshmt/gH5a0VcLM/3TcjwqJhewmEK8pZd7tNPwDky0eKX2w00An4g19
jakehw3FXPp2g8LoRyi5mQS8VzznsXZxq5F5C4I6RKyegmEX9IbvvhN9GVKO2M0HfSrStJNMQSgE
DJmjz3iM4DZHWz8LTJDx7XrK0ZsVt0EkJOOe1PwDXEZOX+wVV/TRgCG0QeNpSFXmueB22s0SJ6aQ
gFi9G+RpoldGfQ4RLCgI2Kjj4DKUks3opjvlQpNpd1ZJO/8YWyMM00Klk48g6L0552i3uiMyef+W
Dsrx+D/Mmp5ivRu+NRd1kC1YNLqb5xafXxym0dgpbEMLrlfq1A8zvko0PlRrGSkGNAdWz87/hGBV
4WCtDOryQQ0VXNovDah2aabNAeoQu1UFlqqgLiB3uRMduLZJNpOCAJgfAmqPK+DJ3A7Qb4lgPGcT
B9naeJa3EjiSCl6JjYxkEq9upJq2ZYI/6GfJVM5bCfP/LEJKZ2dp8ib19/iMG2NEDEgOU80IipKi
r+qIEyiPCiuMVCP5+7zG1+97WBAUGyvUyFkhnuXQbdL3zpE4G1+tD9FMTT8rV53vheytoMoKD2V1
j9MBNc6EMZvHMcMlhVEOdfxZiTD4vWJ0yYLrEjQ3tFG4LTApcMn3HhpjpgrX4bVDoykm0RtMFadM
TvN6hSSuuj1W0TL+3llCQKJ0ZxmIy4oawizgNjIwVnVarLuCOLuD6tFJaV6X58KMWrgm6SBF+vNy
tdBmiBzqYEiC3BDKrXssMG5IHnXXa9o1jVWoFmYpBSFkYTrpFfec/c2SJnAJULoDFobw9fxQ7GNO
zBobGvsiPuzC8WqE+rvgdMNARFQ50i/1A/BlTsN24le3Rt+M1vmNp02JtNAyR42eMPDBSJQxx85p
4Umr/SjyYA/iZ7GQRit+vgNC5AdQ0IlBhpPT7TpABcNPBUxkKMLMEOe1hfvDqtKRUOh2C+hhSZ81
Feu9qLfdmDnGHyTRoS0oF95AMQDI9hBX0aVw4fsFbiXb3Okv75HE8RVFqoMIyQsJw4EoJQTSMez/
gDfuYXh2OFhEqtHbi03phaDoG3plF/ia/LVGrWsHICeAX4hfAbuk8bjBabiBPt4lcfCVn6mHWFDE
WoRj5VoosSZNQsxxyVWwXdm9HGHZrDp8pvSrJIPLofonQPkVWxkVMacV8lQMYmLZ5OjmS90/pxAQ
QGo2lwRKiUeEpduNc2+bZg5r4z5hzaO0xLcWjVmy/V0aKf5wG8WODBlXFH91b6wTlwCxH1kR9GbB
/RR3zsiC/EC3gLS3X5JxTHZIn9qj8ugS4R1BRefj26issatkhdGR9OLU64oA02xrdZQMKd0QzWsO
a5/j5Kl5ITLDTXmJuxQyU4tM49xIa6f3lbBw9sH9tRE1nv/j22RmKJjyVz7YAXaKTFCLbZ+dlOuJ
BB/x21ag7PXzDUxbWO2zbnhagltkWHURgiIV2jhogK0N89arY3E8AxItZltJZv2Dwb3FwDAVgs3i
C5Wri5doJXK7EiQOlzk3duWnOqnkmTUvzSLrGeRTD17MGE2mag6K67hIHKOJQNe+ZA8hgc9fcvga
vrRu4fNKQpiV8f29N8DJlcoGUfoNXwXS8IQAAFzWvaXlPXRZrru9irwS+kZDD++1blpbQL1rF5qm
BRUuyhdlId2ug9t1ncAeLetajNQfxPEOB4sUzgiAU1u+M4LZQ7FM4lLxs5SEuVNK64xPyWcRXnGV
GpFibYd3bHRpsyWYEoHyv4woZNDPFb3msqGcV8fJ4elOnCNHzX2nSa91oNxfOvqO64CS5KkjLCBC
Pvug+rMBAIqkxy06N/7p0VGcaNYDxPWDkrRPhdkon+1mVlpk+yzp71zscBPWizX0X6iNIv0ckpYd
SJkkqRfWv6IaKhZrHQFntRlmkm8GY66FXwjNAwj14ARHcoKPgsri79E3u4dXPpe9UnPlMf5NZMl6
Cwk3fTN9i3aS+vUuZhzZ8tC+pZSIExJL6N6vD4AFfSv0f0rBhn3ucH2KE7BP6SLMPQK8GUWRXGsL
J8o746TNPv4spozuQVnAnY50yysn9U/gsZVED06onzclIW+WakvCpOvXeIlzYTG9XCeLR8q/0Y9L
fdnB5/jB51RS/yiyNVcarc2vxZUNDgGZVX9/muyEUYjHDK/3IwWePc867lFIt6EtpDNkoUvw1NBv
7ewiwUo9LoBDBPYjEd7B7BUhav6OMqjLqnUgQMiGyrB58lIitAItuz0L+a6xcyY4qDmXpv9lysj7
4bIsDhHNgkJGqYrb2tW+obKnH/sq/eOMxfZTmVRPuP6JDrB4VGfWnKRwN37XK2lQMLzKSGr1cw21
ij9nGuIHFPVaEblXsSJO0Yyr/odyaNahECVHIRV4zcqBsU4FOyHyIkSwyDC7fWQ7jGxvYXALmmpO
MPI9M7VEvQOs5UqCixx6diqtF/pMBDt4nT+R4M5tm6QaF4YkLuYZXqsEr1ytz2ycVXfzotYwv+xl
z9ctKK4JS3RgmSPODqcnkHePUSTVM5PKMXvsOOATvx7df/4TdgTf2rzqF0A74wRCiWqGV+9285fZ
Id18r3BR21Ji89lE3bXXx0RBDAYf29cX86byK08h8RYpB+lb1MA4/pwsalCXxC1WQmrGqzG+da5Y
FY180oDwTZ8yRP+JViVu5RGA9Et7XEPERyufoA1H6d4t7OXmJCaf9LQKIJAooyIhd5aJD8Eap2JZ
zKxe8bV3V8cXqVNdBbWzdZ6iqVjwnn3UZJ9SOZ30XQqQG02K4t+hQ+EEVYtoSv/d/z5u8W0GnM2R
Mq7EZt/NMoMX84qCrpPioCvpJtcp7eqamkYEtRNFeVbLfCqCplwm36A1xjfNqLizCEBsbytPeC31
OqCWkPxtcbLuvssxpwNcla9cWOhCAinSTgb4xojsQUdjqIq3iWWph6ajZpMiuTMqWmrnu33YyWnl
QGBTr4SZeHb01PqUNkEgv914TsrjFvEzSOAqsHIz8boTs8OneVJyz2jX5s3DBbR3Do27i4cimflN
EsYH2NXGiQK09NvASm2U0jWCQVHtqtxSgFKULedivGn8gOsRpJk61WJQqTMOLo+RnPNfNP1pglAG
ayyH3QEHwnzdJ19I+PzZCQZSXIzk/aRs90tAsXULGXYBTT4+bTum/lRNuApI2f9I6hwiwGTjnEP5
q0657EKDKA+Kn/uKYieG9byAJQuwpbsmeNZIohha5qWLXlb+HJ1UOWPclLGG+nHqAJ2Yqhfy+Ccx
fmblqphcJUML2mE+rr4vL1lWBqtbRdiUnPu+YxVP5g/jqecQlZ4UYdzcoAaZc0Ie/HhorgR56OoZ
cl8rUk6nI2KTRC2ZcLWXqdAuzz8seZHDf7q30kffoyNUB/eTApU6CChjHbrMtn/Bpe9Ui5Uv97cx
sjoRG2M619+jESeud31b468lhim/OdKx65wGRXm43ktalZ6uVEEQkhggMOjlW7NqRDJdG4gQnQIx
6yQzeTqYj0h7qhmu0OilTkIg94e/9Pi+ZEHEI4ZW4r0zmBzXpvtUuq5LcQ/XnAVWYChcKiBI0wEP
90HYoX+K7l+noYPip8OJYtPNEgAphNGAAWsVSNzPUSC5X7KyTFwjju3gQ1aOxv3UuS11+YA6pfsP
eNad/rOqHkHU6uxiLF768vN/Ej5dQ3N0B1mlRPOiA0/RMfDViR/4nKQKSafa6yiIay/bBFWXteBT
wEKSkYBHBXrBAK0BMqYNYps7qu7Ga8+I7fNyRWT7FFNGQKfYvYXn1mGT+rKH40boJlMzyButp91m
c9BKI8+GiSNBVoGqlFS0bf/9CEURo9gHigStpu56SL0It0GE9pUjkmOsGL4ZIdc4c3X+3jCDO4xL
Jg5+eQBRxe+8czrn4LAlx95c+lFmnG35rKZG8TPszFcSLFf4FxiwKHkU2tMN1UMyt6muEwH3DG8t
5hD86Ess2YDkYtXT0tOHkBt609tczico7/DRityOJHYsdSREpq6DnW9ii2G8XCkT1sagFc8fzMrE
nkaYu53u41xBdW3lAz4NZ86sjig5fhkRGsI7IXZH6cFTgRRxtmTaJuICGNCpv2g58+oWFO05T0ay
XeQtxX20YoL4cer/zIaE/HPxjpx/WAmXjyaqKIZpDKCowIOYjMyxqo5nbQWtUwUMrUS/SiIOGEap
fsCG5bB2yjuYmsNwnO7/px8xim+BqnaFe4AXe6C41HLab7BbhDxZDZcBX+ekCWht+zTN0QIOiVW8
1+ieeUrOfCjFOy7MqyCIjMO3us4+AxNvCOnoZUlqiMKQnsiNe13rxtOkVFOctlIxSX0x4gRhN2RI
P95EOnwzfCJvpdIDKGSli33x4wZYGX2xTJurHWl2hF6fnnRAWxUb8hNhZiQ5n9MjpiC1rDLFRVZq
IIgHcobVeuVSHW5+fYtudF1Fj73m4Uz17bV3FOp/jhQ+JwBlIm+VKRuVZK2VF3nCObPo2Rh8inlU
1BQS7YUfBSxvA4FI1fkvGINq5YTyTVUIzICDs0Sybj27kcKrJORE5+JZoSoThwhJORCR6RmatVsS
xzBo88oN7D18qDMU+VuX2OZp1754Ymu4JlXuStTbnuXcjkPzDbUI3vF9qm4T1qFmEp1Bk88gcLMc
kt69rSWI4cb2foFniBv5lbcpKXs4hOzkPZsUGpqAZR35oqhn1UlgvzBoreRRJcbvFjrAe2t+9IIE
A0Fbjni79sH4Rh7ulamPFIkIrdgnZDe65UbSFdgC6/R4jC2WADL5dgu66R3UlAFm4M6/ys2LJu0u
xI9kEfP2FcyDwkaUikdfhw35bVWXbKZIpdEfKmq4pn2oO9eYQ2ZktQuhDjk3wYvWvFu8Qd2Rjopd
SrfNs9vN/Mz84nBIKuu9bGW+dZ55IZWp+xKY2/vxYUb9m9jSSSG5FpgLJwnKkBY7NtkWMlHpHui1
oOulO1nlkrhFHGDFgWaH5GiM9YcZ89SUpqSHvgOn3yYZMOCMBGy1K2gRVOtOUAQyxg/1WVxJzlJz
mAk6Ap39ZLvAunoFrlA7BblWDflx0TcJj8vM9oVvgIhBfVpkBR5OkTcavMlukhFnhaholHHOa1de
mYy/neqWgfkJ7Pas7GKc9BIPEB7yEGBVkDCxleNPXpA7WP0V8GvXZ432c/qUQMwWvOTLF14KXHpi
lmggKoyqnFcjsvfyVQNrK+y6b4fyVT1BjA83JOCayKy5M6NJc+H4mRkki4iE8ZHY3ZV5EMOpWWk0
aMeQtupbNF3kKIeDAyx4M6R8XRbKC6abw1pdMCSlURnGRCXRUjnQfYAnd3+Wyh0VhH2P/lNBtNk4
cvapDobwAfmueijLnkM/mCJhshacgw1wlsLFc3lgbVhlUdCSGIYsnp/N+L0maBA5n+01ivgP7+Qc
HLvpIM3NLa5VWECtDPGHVjbq8hVgRq3EAua0znB6XIw3m1WbwfnELPMYQ7OHPVfimqPlC1oAD+6H
mqYFOgELLM05Hh9/Yce2DpLoW1CBFZseT73V+HEkeyf5hEpOZYEffmEJa9yAuKXos1IBHPDP/jKa
1Xju2aI0nsfzDj0wVWm5nh9fywu4hmcFuiHAE6qSlx8w+8yczefWgXk1BEtPPrad24sTqsyCgtpG
bTH4xg6nz1yKUlc8nna5wm97YtZf0a4o7JSoSRlPX3vQn8WnnXoim20qxetU58xJxZbUFlWE7VoG
0pRwoIsG8hDRZJN7KdAs/8whZnhph4bMLMcaHPifPic4/i2pqD6gUieReFD8j8eee9U6Mj3OJDsU
rYuCkRW7CyAnzu2TZdEmglrnnQhmqwYfaTs9kA2fWCws6QKhnoTN9HYqqJ3/W2piYX/okj4xapjz
69ANgYnYnUdmhZQQliY9ZN0iQDi4T6It9f2A0602P3G86AZBrP/qzvupGZ+8C75eYRswxjjKvK7B
XvSuv0FYXpJ8La4EauLZIhX3SHSYVgv7sV4OOo02/RGCLNV74KftY1IkgrNhZHM72E1Vva732UVB
tc+jG5kKpPNmeGhcQ758JWVKdgyJurt4D9dRtpH839scYCWJOfLyBGh+INb16TU8cRVg4qa4/8cN
/i6QdcrYiNTFOG3mOtHFunep9Ut+6NbTiFYnvbNpRCdkCiRf7YgxgFy2IgH4j2rzAXqujcwwo2JQ
F85xwt60DMEHxqMeHbJ6bbYdP6T8mSR58MLrLTOvsrh9Ye1V4o/Ku9BZCHsqeUrE9veKUzDwB+Ms
DHUZR1WsCXheEBAbG26r1G65gtOpc0XecogYd8ehAy0b00fd7Vokg9W+ZxZYQT9etJ5y+fFc4M5X
69+X8pJifpC4BeM2c2/CcVsmTiyOdQgHEJm4V3LVwSX7lI0rwd0NYAzzL65xysbxvQKjF1sRLnlE
CW7TjUV4ILCbC7CpyNlRJQYsdbSgCVSxN6/hqd1ywCZbLTorbi08rHZRM9IWLXwhVBhvOnHjmg+i
Ig7HlGX1L3Ow3ZIR94plPmxeXrazDzkyJ10UIKuDFP7U/62gQ2GWIaLizPSI+zRss6qV8a4SL/1i
k2toEH5rIbvyMWDFCavKIiiiU3hVJlpWgd0JqfTHD76/FAL/YfaK47HlJCMbHASHmh71LO5v+gwd
4Q3Gna024qg7CEBnlxVpoiysiQqjRyGgAADBHIQIiY3lFFDYJk/Zvx2ym3GZfKLZLGAoRIpf1X9b
7sINUWggG0QoO2xFIlTI3XHl17vIzi3gK5ElnjXKiNrP4a9DEK4E5fTA/CbvWAkoz7EO52Ywi9E0
z0scEkqjf0NI+PYa9WH6B7CGLGgohQPK034tVfZqGZz79FP7f+G3C0NqOyQgSHzKIRn8IUsNXQq8
tmVYYP2fzsstZumirxJp22eGbkZMA4W1YUtWsZ/8U2P3alOBfLb20v0HtxBNyVIiEfZuFMt2opEn
Ayz0m2azNA9nmpIhlG26yhY2lUKzT730ySHoQDA+aUm4MoqVt0OMmApqNv+DNXquodszLhUqXo2a
bDIZ4aY0ZhqMho/aHmesrgsVumD4fb6FYqx1d4t91OEnOoogaiGpfpzoQs8d9MXhyBoQXWyIVbRy
wHsl3HICcPYxGqtQNlWF8XkZ2OYW8Eld4ulZlaHzy2bfYtaXgTwji69Le+4qUchuUjICbHiyr+vQ
P1fnQaOuYQlNeWqUwTDc0F8N2aZ3gQLx/X+LRILi9IfW0amJ9zFvKO3kfXE2wDtOadvTZD9d3h8F
ZDLwpL3QWJUWZs1vbATIK2WyGVxJ6r9wKawFV/7zY7dR8zZQDjlg4dF7oCiWrneC8MTmm5Hd3Pbf
VkvfZBaCQZD0N/f4wU0QqpGsOg1uTE0WrvttQg02VZudszuGewRKDYuX5zeKVcHqabh8Pv1c8hQK
i06Nqg+RQZOAXs/UFw6i47l+5iEu7Fw+qcoNtInkx/CA/I6lqJpcc5ftrRRH7HbOUDT0Bi5UJDI5
fIKhEi1qiHsZzOZO/YTjZG4iM3RKyqKMvSvKAZTv1JmF9CrRIaviGuvG0+UJwL0RGw6MYvSz3Uu6
EgX/0EflBZxaNk9E8973W81ZtMZE6gqMyyAy5QBOvbg/b1l73w7BJg6AbG6XMjwa6GPPSZiEjMO5
sJvBmzJFN2gZvsRwzh4K0SsrgYn2L3FWY1c40uOvp0Djvyr4cUfVUDarWN91SW40lc/xIfI+FX+G
xBaJHj4OWXVog+9tEZca6QUORIVocpCPiAg3xsDIlHgnndKTMT3Naam4BjvCBd3xhEwArr6FFoOP
Yv5jB89/kwyXDqh3S9N7R9YqEoOqHkJGgJTQ749hf+GZr7u8zWQHEV1bYYjTgyx2vqPTUD/x0RNV
B3lHlxvXxgaM6Mn35Ve7qdg3qoJcyTjNt07o+k4G/FwT9KfLUdiHgyeBPoKJygdibiL6LN3XDIe0
dcwWIiQ/AfuzmKvjY/MJCrTLzBZ1d5+gOGOua6vSgn2FU08nj7X4x8QV3HdSPoyzCQnhjD5+e2VS
zva8kWylLDnYGbZ4eRsENA4fnYvzyHg/bezUhhx4QBDDzjqvj3dwcwlp2SSS4fs8reJhMKW8hmLP
vbCSbuDqKFejlNwOf9MOkiSsaI9wzcf3ZqOyrHqmMX6xHAZXDQR54AmPa74+kjBskMZ2OxJdDmuI
FzVULF/7YV1UcZEnZQBiP8eEqB3zo54xU8bbuQygNIKcGSYBUXVnRw7UXVRlMO8Lkv77PyEHck7K
JxtEG1FAVm6BbhSVLk5+c9MLM5rD7Ww+gUQRWmdcidVhcdLVxzIGMyQ5FbeUp7rz/zJKF5jQhrsg
uxKo0yt4S1r0VX6v+a28yzRnsH+HP8HB7WeBRU0kpi0TadEn0J1ktNBd70mGJiQehdGer6iWWkA7
Wtii7ERCQPPTtq7oJYwXs8t2PKwYtXfKoUQNEZ4SrLiG/BJtJg57ROA9bs/WO2rti87bcqxQQPIg
ub/DSBYwc+ORAjHjQyKxwQ2L8DkmsRgNfC/85HGEDCUTFrFue7rWmBKuiUtuHg2VTE3XONc03AVZ
X86QpD3IgBiYk/yyIhdK3glSuh06N3FbKnbcByTIgR3kmNapopUucsa5ra2Oc4fs7esSYM6Paw8P
S2jG4TrkiAD9TSFcdCtFW7nxf6G3q5vn0n1kCzTmC0ybo68fg00oAVRVl23sLEMdVTOG/NC1Klwb
ak8NcijgJdR6Lqrdc6UIWdl0hwbgX6xaQeYRN6mqlrO0j9/RPQQmmF7dwRS8TocUW1Li4qV9rbjJ
tbhX8hUg+SmuDjXphtyDTS3nRUo7QPX8CzpQK/lHfKwVxuvUVEFBq7Ro4mnwImlmGGJXjFQDklyx
J2Lqeg3kOIu/AMuJh5TnvaM/HLWCjsFgiQEAZu4sgrFeZ57W7Y0Qs7H+R1lpOE/kb4oNdOWe0fhI
T8xF0zPpMAQUk4JW6Q76ZSblk/roGbL053Ht9VLk6KQxP1D//FvFSqmgIWLmjj441ROwEygjdqOL
pYoSCwaVU+j/3FePJLL6ZwBpBvXfllCRhR7el6tdXD0Lsp3B1ZbXrbHkQZhLCSP2T9Mv6saXzKQ+
lszKm7VYvbnMhcVNwNePsHkZTFcMC+UHZM0IJsup27ajrUGs5Z341wVUSSgrHPZLrDjwdKJN6EyT
CbsTRPWYzhnHHSm2W1cu7girJF/phslkSeTKQd3ax0rFISGKCBpeGZopHFvc83w/dI7FwHb1ySdW
pv7fYwFIZeXjehDnlGeTXSY3WBgCmKWszSCIC5pa1TxOvfVNOtd9dqCfMTjUaozjcaYRF2Lz/4WT
3JDuo3LXIKw9Ijt4znP34Gz4oyTTPi5fxsDDiD2EhUrmdsDGGvQddwmmLKqcVkAS9m92W4CwTvjw
gim5a+/0NVQigZ20VmVy1y9OEjwDfbMCcjUfpKZjffEREIqIdXi8Vux+VVVHnW/bNnTYm34AOPZT
VoCFMefb/ZwrCYQvZKXuwcr/DZ4WCaSLekH2ACNcvTEV8EUTNpMFL2YRuiZxMwEWA97VPZ0TfIZr
Z/pQslUEzPwOz0lF1AVMgPGJindHR9/+9ukPKSCOdNOTKw6HHopg2Bv3ohp5PjOJ+bcK/WArHETc
ShAKElhdxTRILW4GqnJh8U/Sv/h2bC/qp+x9dexS8LxUN56VW3zkklzgu1VdVGdyTigaIWEPw2ce
bhEp8DXLW2uP3W3Xo/THnS+jrTU9Y8FcrzZcL/GAkchfcHAj4PIIw8QatQ3YdK0Vqw1Tm/5zC3wL
QipQf+VUoPUBgXfS64hwEmfZtJt7z1Vko3tMvekivvomvkOC2OGnBvq3rnrP9EWkMdYnaeif3MOD
i+XGOkn9Z8Uxfo/6wc76pnBEFfiOuXDx0tFLacyPAw3Nuw6ys9N2dgFD9jl5R3Q8+MLgxxFAIrWk
TCxwnwv8JFjm1d8e76r214RP1rg4aQSd0RoGWyUj0aWok5m+bEopcMIwG2CPMh+kXUKtsetGlLas
3due61OrXdKI5At6QTdyM73f9Vovuwn1Yy7eRvHDGoYsi19a/ZBX4Bj7wMDrrl2DEU7KLoAAkX5y
8/eYMQIp0/ylhkjeWKiOG+bqA/mKVVWzbQEuzlqzH1o2C/lbmm8p26f66ab90KplWLO21bMGoR5a
hYZj8688kaFF0v3J3qqs4hDhWSUt7zURFTa/pcOGWPQFnD4DmL9PA81AxXI9xyJMB3oKALQFqjix
Gk2Yv/pMNbstIHw34UNYVOtFo4d6AiFPDJRe9pTFc5s0JVbtiQ2b5STfRvTS0DhEfrf6/zCZGuIn
dgjcfy8b6mHm3wT3hnXTvdb95QTSNgN6gKX7/DQnTrOwoWjFk7K2ea6b6RKtvO6fjimNkt3KnqoF
cbG4IrCYTmiFaJYfUU6yjYGL2iqizIQhTIrfyeeOBqQb09LXEhT7Y0xofEV71kVWWkUfx2D73hT8
lxBeMSe+laebrMeNQBp3sAop2qPoclzPvPyGhP/ozrGNWEM2TB9yU2jW2vYSLZwvIFUszcBBcjsl
mcw98t4/t3R79KU76jx5AMgvOiZxa3zcEieALD8P2nx+ENdfvjYg1d1kxjDGY+8DPvfjkAasrQPP
zu0Di6ep7G4YQlees//b1EaYqPhvCtngZmiqmNYYstJQpTuE7iaPfq+N5iu8h8kL5k/LSSmxuQx1
/zfsY9OgRxXytC5+8uDvAvJW/i18pCHku11+05eCavjCuh6TCrsKeFgL/OTnx6sMFJzdYbFs5wxv
VYhgTvz61xZgt20GCU0tsb38GNhdPATXy1bSE7cQB/1+f92zZ+S+cn4kfAg2Ap+w54bH95qi7vqu
KiaTE1LgyIyauxmQcK7RVJx0rBdLvd61Z7qC/U8kOC2v9uz0F52q+URJqnOMmjLNGowPNEf5uDkY
0FNJBxK1qx25IJEQsnydknxaP2/1n1EBKca0SZStch5w9Z71oQiG+o5gUqL9DqeWuqcRMbNpxi8v
auEhFp+gv1K09ViTByDK0Pon/KTfRuMCOxtvVSswt+CNiSo98cr3vpYbnGxhWiUgJIaYnjdogDXi
z1NXcyD5z5BWaq961QRajjCAkEZMCFgQss7cCtFz3qrXUh6hIS/agQulCuoaWAENsNMHGmWDpByq
sE3g/Vytp+ou0DySGmDTC+vV+Yi3xkF2BVaU0dc3M7wHSu7L1pqE0QRlGrzIR1HBolZTL51LACjd
aDFZ/t2hT1tqwPiwMRJnqGnDjZhYQN4ieLYxXalzWsiGgV0kt2NJ9Oba9UKeA2DkAPSVTHBAa1FF
T6+Ft4rhHOglGuRXu28jpFKRJkYj5yFPeX0cLifJ99RrhI9l2rSL4b/yLa7BJdI/cWQ9VyUFjIa+
ci7bVyeOUgJMFE0kEWjbD+I9V05a5WXWc61/eJW7EiHrJVU/x+Gf7Choox9U439T75XuVc1GjtHv
Q8BO4XDZtvWwWPnjWnbO13uItuqfiCT92PwwrNR/+fLcvbYddP4HGK/OyHRHAphBJv26Ta9wkLR+
/hs88OWJdRwXA0X5tGARPnyR7w83wInPgU14B10P7rYYPaKnvyZWFFNZ5r1ayuk50gYsim5+3O+U
MpnfdLaugQhYnzSaBMK2W8JRpXSqm9QRw3nts2ubOnnwtDejVHSIu0PEi3V35apsF3sFOdDs6Uo1
ms3+nqe444bO24KI6iM03tQ540wK/IpOuXZ/g9k3NUa85SSBDo/OdM6Vg5GbtMMZAmnj6FY69mbl
31r9PC7KwLJs5B7rrPVoT8KjwLgH78XINHiv1TUKuAxadh/qDw2G2UzocrS1Li8XrICDF7Yr7gft
rF7PO1OQ2gZ/i6NFOl23VZlK855cfAsgHttznruPouYUEcWdPYst4uDxfQG/lPlm0+nGsapvrSN0
0QiO6HKrucmaTqCyfh6xO4LqY1ivbMRimA+ecbVEt2y/TdWZE2ooWUi/q1FcNQLB1fioWZ3qS4pN
tk1azdg0m5T5VCDESXYf2PQs2BoXfJwRmvMYJSEY0HQUdhLHHaqshQuHebR5bbHDBg5tIlbh1zye
4g75HxwTCj4HGb1mPAMJjvMiQj1Gmx80/iEI4LQQoihv78AC3dnvGBvLov4N61CrPZdkL2EQnBVP
S/UR4J+OVAhIdXs5KQY+IKaJXZvmEAjqQamXyv+ZvWVDOZR+oj9T9zamFNUddfcyROrmcH0QrpuT
A4YCB2+KhV1fKsiCZ9uS9TbtmNjlSAG1DJCfw2BXXwYGFCjlnBE5GGzpqyW5dCcki8x1F8enbqRl
HCYluBctIVbAlGKUoLeY6/OpriN2J2IRzswp0wHRFPTeCvjBVOG7i2cuDej1KM+7X+HflGrXsn1q
o/iaT9iXB/ncTIYXN1NDylpTySI3zikQG3ntiyai0ye2g/gALklznF2Xw7q88hgW7gzxh8gueEbE
eh74XYcT4LQxm+EqrnlQ1ZeZ8pIJK812GUhbvaPUELYT178AjUJ3Ax9ygCC9fF5Z4Rglda/V7E1r
tHMoi1Z+wmrLRkWONMsvULkC6hupFcozwAq7rdZFPDMQYMybY7S3nqtCKXp4cwcoJejXUXgjX1y+
lNEgLSc+IN9LIY1Q1ZV1K23RXs/H86iVraV5reIfKSC2740h+ptZ4CWyGQ6hA13dvZn+iS2euSMB
gOJUBMH3GF2j0eiUVG0LsDHqwQ5RZVamkaF/4twIGkR2Z0oWmCQ3Kpj0nv2UjC4UkGCWYd7YqANe
ffY0/fWxkRF4tI+ciY6V0h0eJ6Q1cMaYHuzliKZfQpAUYX8ZRbKGhMCCIt/1FWSB95+oFU2A0N22
+kteheboPaQajUMtzgFdSNtfLzs+jSWFFXOh5n59QQMIxuwb7ydk6A5+3e6FsOv6fT24i/pQD1Ta
CZyze0v9x/l518DJZNXzawAKsRnAKAnOnF8u1swiSFwil49kwPD/mW63Hkmz/j1zpLXogxz8QDLa
UB7KyvysB5QI3+5x8VzkaGAcamoyduy6yFIqtV+sTUHasFxUegr57AH8/aMXhcL0Gpm5lhSQrNrr
aUtj8vlOGswvRPJUu6DsKVhYlJseMAz4zhTEaRynjRtlyxfUeEg2rnk/AHulAcvSzFY88m27NbSR
nlAifqVUt8XuGaWABsdpl+vbMxemGWz943z12Fdc36MxF4FxYkEi2lRwGZFHmDcx0dc2sdHXiQm8
M6Mvqq+QY1+bU9lIGS08zt/36S4yhaMVNrxEMllziP+NpE5ZkMsQxW6saP+3sYCiIP9K9P9Y4TPC
FuY2BQUkchz2C5QbMx4bvD++82ELXrSsvwwbfKXFbDied8elYSU5yFcaQlneIgtK9LES20uAGRP0
kQLyyL5koX/offmAzTuuTNO+2NNnXo+uDKbkYnhWOSDBjYhnJhGlThGHRzUUvIjAMOKKCyqlFSFp
lGL80Z74sjlYOhXUD//Xx5lRVsbr+U4CEhKo0+9WNWQ5duVdrc97u3IBZw/T3hmOeP2nMZ5C2t0/
XSt5fKnvZyLtAB9ZOSdNjSWzLZlTX29Ns3c7VPiqJrxiyzsz660ukddEqjBVyxXFBNZeXXreSZwP
MyHUC4vp0i2JYgX4PBZal9IzBPaEShVnZq6AqIVnc+K2AZUq48OE72LkCBPHfqeROQzNRQSNxF3Y
DtESKz3SsqxlbKmVPJJUJJ1ACazVCRs1gGAqGKRgiHs5YQJI+c17PoUxthD/VQfey7HbCZHiWQmy
BFY4A5XXGl8b+3t8mHL18YFgoSznvnjEAqZeb70o/+xRzH2KDiNtm19YVlxtrq4Sd/XhYOSZmwV+
kEoZjJf9G46jsSLZCeS1FrYHAqVXKOykeValpD8wi7k/zN9RqRWPHgvc4tKHsxHJ3YoaUS5Rv6Rp
ieFujqgoYStIyzScCB+dAWTlW9RsgKXBqlXxb8ydUQ4Pu5RlXhVvGzP/dgJPN2+vV/ySznXwpCe+
1jj4zzTDzBvAStL2qGG2RMhq+AN7D1hrA07ogLfuCpNNj/t+mwxbCRoSXcFVDnA1joG/pV4pm2ED
m9JStC5Q331HZds49IAi7Qqhap4NuHFFTlyffXO3W++jpO2cTNRE/PSLk2V9DB9Rc0SQepvgIz6b
O1j8KJwyYBEw+8ab31fJxmwrYimAZiy3aiSwo2em2/r5kHgRTreuJWlp5ev/fec62VqHK20zAHIX
TDqRh28+Gm/NOcAuEdrkyNX5VUcO9lwRRi0UvBu7XrzR4pNMffs58KWIT/Vzw0MKPvjJmRihIIys
7ti1LCpKuXz+NTsO25LScuyHMStc0TK/aSQGGAogO+ruFAXm7Jxcfi9a7OU9t7G0Pi5jGJRUy7q5
pbbC/kIsKKMw26f2u4kOJMWBSzE7QNhtLq6xp7DkA5t3DW6n9W97mtKp+4u7jYQ0cjdd9mtTEuP1
TB+66rHj0mZXHaURtKoTv3Q8L5PGCFHUo0hhzCRVEKVrqI27BNsA6Gs7K+daSyFx3hMCsCK+pkrH
ooB3f11GjPxKwXO3UTTwa6LrzPXgpN10wNuBdV4hu1zlZEkwQx/+R4Wx8yZtcC1UT3wKTOzTfFFv
et5xnVI7aVEuo0EcJeRAnLHF7KUwdSc+jaQ6DI3knFFM98nEV+XGSx9Z/vWWMUhnACDFcOmiubh7
X7qu6u6RdOAY2/76bNeObsT7cdKz1p9K2evFEvZaDUL4s+xHfrmc3684ITIn2j2ZbCrvA6KjNOnZ
vsFDWVV4nxULF9XY8GVUqtRqWamyKRzkDkhrfVaIa3Kda5qgNPfAmE1Ml82y6XGcN0ZAIo25XLJg
OgOtQwMSBOaoHd9LTtQ93nB/BS5XHotQV3ClOT3ys4U0MkTqzR6G7uTOVj5R8r0GT0V+P3FYt445
/b8+glYfK2L6hfIx2wYDBhWGz6bWIcBCrz9zervAeDtf2W0t+pr8rQLgSrNNluJxDc2sd+BVVElD
aoZjGe6nxjf0vFPBbAGW/qQtPGimedWKZqk9hrhqvu88tvga2wHI/Tdvtv5oIahFU5rMym5Axh5V
F6MeOOHOEB6SWUgg5H9WFfe6ZwFD+CuvgmOCUgN7oWqKM98k8R56U49SdfFUBJ6gYPRU21Hmpqlk
ZOw4UjtXuxMiGx9I3Ajlk3k7CFqjXN1zEJLq1HwfjWbhJHL/zVCUYAMor28zIvRRgtAgI9ryrDB0
g+N2sU4/TrTHGIQw3Vp8LIh8vnt0wEvZrnyf8KBRfEUwAFcIS/W/TL2LOPoGwtttP6XIiBLx4EDU
wFx2oSJvESfTq4Oesn2GbUh2Lb/SzfE/ZQIvICQh0wzKVSHS5kalPxXyWLqhi1PZM+Qf1+u9c0SV
H9A5oGjDYnub0IvBVZ19/p09jsPRAwJuq1ZoYEkg4sDTz+XRvKaWeH8GhTrerZimP+agFrRZNRP2
UbaYlYCl9kW4nyhFjY60HlQ4vGSRrcueFUdqvWGRQ7iNjAndHDrix4fK8DhLSDQjp1pvdXFkqAp9
k2sVzUBxmNX6igGxSOGHwSudFLwOkMclLO9QWcaassFskb3lExrgAoqN69vSuasrbvg8ALLKj7q+
wzqnUoE41q59ADL05hEwFsl0VTogepucPlLu83OH2Zj4+TMEeghBIo9/FeB0UPK+Wn/Hr4ecPmmd
bxmaUkZveniZBIVJQlErBVmC5SMd/+aFhoJK7TYrz7k4Kp4rAXZXzE5D+xwCD8Uhu4jvNJfrAan5
tPgacEP+RvQITyZMV09Q4ZT7o0t227RswaHJzDQDvz5hr7Cxa2j9cmyVjMGE8NGl4DBUYMW4SyeA
/51PB4aHLfLSo2pnzEHzGBYYLje93F71gefcZvdBOeDDIIInrEybFR77j5BUuKagOlQDQ6nn4Eih
zTQzl6Cb45LcPoXeKNfQ1lIbdjnwT3I0EJCPT+lYnc+fTv5fj2kfgRb4hBlIhphmSeQZgI8SG3J5
ev68AFW+IXhb1Q7GDoe6gb33Zoo4rf7WTL0oBi1S79T8p6zlMQKeP2QeLjWaKnBNCez10os7GUqi
oNrFt3H1A9c1XLTeDi14wIIxPW+EFmefiqiWaAPCJmB6sJNI6I8p9tA0PxGZD6MsQAVEbQIl2T8s
RcPpQIqqSBbHnreDVKAffejO0X7aYbTThYaUiaEPB9fziy/Ho8EfWsaqKSweQdWi2Exd/MRm97MV
RPXg5qLFLE3j1Vojhh8MOM8yQluhCni3WhgpsAK71WQ07U/G1pP4sNd92+ImzQRpUVPGBzTaiy9Q
Hf64vOCDvn4aTTgWyqtb32g0tW1JOXOwJGp+jhD544q7nbK2g0Zt4fr0Jkt/jFPWX3NsIJGQWWWj
asSKf5X/4ZONqg100D77z7sgH+5qhrT0R55cC+xPrhZuPMEAxiOYf88R/1w4PXQXY5wE4YA4tdLv
12bhhYe0R0SzsVO0Uz+p2CXqOn+ZlV2d7Wl/boyTwnlOFy+L2ZaZBgpfzVBNV8Px73O6pLHEJN/e
4cwvB3xZdBycL4xa7fCftisvo1n2hz5E7+zDFTZD+VDOTyiWAIlXjq/2EYUP5HpuM2zeT5VpyIca
R0fIpcr52ZJ+sCKO68g3RpZK4/T8Pwll8qQM+J8d5DsiaV4oYEdW7/ATZnm8BubceUoOkSy0HJqU
hM0gBBGZlKlSAuS8NpcB5bxUrynekvSxzJ4XNROzuQBOLJ20D3M/XnGQYbE/vTWpOFiUPuy3/c81
ZSK1MRtp5rHRpoaH65xW50/rYChQI4BY3ZaySOtNBHCBh/sNGGukNswKWko4ttHd5Zbu/pBk6ND7
AyR4TSJqn4KZ1E/oqZuVWXuPUEUNhggnib9ukjtRBFHYuKKsJdJSitLAmTlgmSb91Rhcl3qs9NA2
oP41t5RLLoAnEjA6cX0DN+nDAijxNxQziYBRsuQpVsLa5vGVthm+w3DGwylJQnGqXjp4UgP2rNIX
G9v82amRS2eFrshdyOtlHCucMXfaCIv6yR4idplHqeBV5MH4pkaYHFCfAK5U1CQmO6d1Dr4VJ4S+
vPy1TDx2fRufKmgAKEUqTa00HW0LqdJaLRsw4g9NXMbXvQncPyWjq91Kgri1c2Mb5zUXh/sx84fu
FMpnl4lK+eDyDnKheSLS+oRLFoWBEH5q/00suR0OUW4kDE/fGcK19csp3BDLKfswYG4MtRdqCT2M
CdlMkRtIPTc1524h9iSiUtWeMJ0q5T4qtWsjku4LawTV6hLyKOExcTD99/lUjnTWqr3Ub/CEJOtR
cTaSFNZ8kU5zquDIeZdwfnlePb9LGv8jD+LkUwOjaSDCCAKUQKoOUb3Udcul7dpYnU7bZ/9r5dr9
b4n7RverFUBHJUXR069ZFf+Uz24/IEUUjC+dPirlncnNapB+LTOHIatxTF4I+ORlWxDhQUuYCsxy
xqCnmISECtao6PY5uquBE+Jdzn9+HElWNtzh8/3D7Bv1qUhELzq8xWnjcAph2pYawiG82EY4Mvn2
kg4gYOT/OM+Uwe88+9nCLTm54PkKoNoPkyd7eL2I8JQxBqs/G/OE03n2xUiv1buxoFkk6m0sx6Gv
5/Hs4+fgvWkoUD/qHBRl1q32HS1jRYGkCW6sHp30ss1rxbzuXcY0kIlMApK3NBg+XTwnzn4Lq2Kv
QgjDqXv9LiIDM8x0R5tjMZqcSxrYiblFXN3+bWLe5hNGyhjrhK4ox3jMRqZsavBdKeaDCuzNzY8x
Qv2cZ5EzgHzBeIhAO4NOiGIejU61nsODy+Jkc2rjvXzWuyaSZUGChILIl61qJlncrWyPcksORE2p
Pye/O3iZozpygjYnN09pS53SBrH2Oqspc/WJ8yOid3SFz83LDZgoi/Q52niuK4HlCQlhcgdeH3RQ
yD8qFLvtreG8aDJT7XXDZl9kmZTwwJ3c5AUxW5HgIg8muc+aqepdH4nae5hn1gJ3fnFu+zHDAOES
iWy1vQ6Gj0hhlpI+sxQcDL9xuJJFqeeQ3tnPMUGTigG6TlnPB6ZjGnmxbg9bAi3uDYnXYt/hpqFR
Q6kBVMzbIyoWEmuXVoBWpTiyvHoOqkEpvuB6/BP9UpUOKV6HJ8+o0N06lHiKIp4KdLMpAE40KvHW
3Bs6z+7rR9kJzY5d6B2K2iPQaFYvnoRzj7cYHUcGeN06Vy0GsedSaF4rKL3F5Bh79foKdIb/H9Rt
HpEuy+4rz3fyja3nrFBHDS0ILrEM0Og9kbLq+W38LkCgsVOhNKUMYD5ymoKHkcVqQaz8xnwVLwPD
EX/16pu8bMQQ/xnmAew0FpZ/4Wo8sChxo7mGg+O7yqGVQW2wbKvvJvFIVRmDZEuNVIs2dyGnh/gH
F1OaJBEmZC2bVqGimmD8lYo7pit3wuvpqQDs03ipet+tq82X95NK0XOnqFDlumcD0XAzTa7FPhWZ
uOpsdZtAKsfKf41YsM1YFqVbqn0wn52aHJ5t6qdDc5iRHEVz19LM3Gi+JoCfjXAuWShaM61lJlTu
a8DaffhyU4Xc2v3Zl5Y0HFIHb9x6g3TvCbMWJrMQyT2dmDpohPCuSRtDm7XQIZYQ7IPGGzYyWqn6
kptaWclT3jQ5VakKVv8LdikfN8fDn+7Q7Dz9rKhhFo4scR/1tXMKHECqxOugWoUuv3m2cPfiO4BK
g2ekzMhDVC1H4U8IVyfxtvnMc5AKtxOtELVDlO77zfdl+yRSRfpdPO5kbo2/DI5hgwGlnVIVM9+v
Iy2mG5M4g4Oy20mi8awy2abTvfW8iQHwaJyXlkn8qYb8bK5pc7JRYnZ3yxVWsoNDxrEQ/U9LRRjE
lalXmilLDy0GfK1edqxfhIc04vlxbgO21vzFvFi8DKXhcDq5LpUWH/wpmp62Q2dOlOi/tpLiu6QK
IH0/TW8KRKKvXsJAHrNjOkbjscJEAIszDFV/sTcRpgl+X1zB8COea8O5HD6qxOtkwf0ykbmE8D3x
slxwTZ40G+ohND3n+eL/q7KtvIdj/9uT8oC43TClR/DhTrb/Du7umGEpbDzgNqIF7UvwAk0SqF5Y
8XudGTIfRgff5EmB92lAT46hXwObrfg1+FLGCyJm1hk9EzohFZXjpD1nmrTWIahwl2+wqN/bJRSN
xoBHfvf5ajlL57Kk01I0jyMIhCtAGV8sqGVD/dKushN40AWe98B8S47msvwHqpG5B8SM0petosiB
81kTT0TCyqZg1ilOeM76qpzncRUOgEYT6WOEUC+U8zdyDHa3+2cL6WnOchSPehgaBsu6PSAdrEaX
/K5YYFZV2LEcjimdTs80LuRynmT3q7qoYv1ilWCxbenscip+vr1tO6R8qKYZqO88l1yB80t1sj3Y
+3yLEK00IhAOTCRyAyo8FcVuMvA3SBFP7f9IZGuU1WVlCGEQiGD/MZL8n3msR3TuaKbZUI6LqC6l
/Ax47i/gbp1r69tVWptsRLs3PkQGkI51Lx2SLohlZCbcsYpQpq8wpOptsTSZlGuaJzy2FgbbUpyX
spuZt3ZttR1iYGIAvqu8XAaLs8/G3YMC+wDooDGbtiQhmtQ2DDmWaXpiX6nJIUM3bdXWVumg6zO3
xRmjJsNLqXlBn4Jt+uDcBy4UUD1B5jzGyjKo2N57NEN6l6XzBkpQSw0vaR9eVUXWBbLl2tCVx/2y
s9vR1K+BWADXS+k2uVpTw6EHKeSggWxsATvSkTMdne2y2wiQRsHbe9r7hfpRyRwOb8NpXYYQjRFa
Gxfq6pyg/lnbMqKVOuD3gFFg1vR4oEdqnGCkdj98dT4Q+YOpvcvI6x2g+EhOpIFYxsDiWTz4ZHHw
MMPW0a8MeMVrP5GvgBVvyrm6OY5vZC8s5f0Tow==
`protect end_protected
