// Copyright (C) 2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, the Intel Quartus Prime License Agreement, the Intel
// MegaCore Function License Agreement, or other applicable 
// license agreement, including, without limitation, that your
// use is for the sole purpose of simulating designs for use 
// exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
// ALTERA_TIMESTAMP:Tue Oct 25 01:51:03 PDT 2016
// encrypted_file_type : local_encrypted
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent = "Model Technology", encrypt_agent_info = "6.6e"
`pragma protect author = "Altera"
`pragma protect data_method = "aes128-cbc"
`pragma protect key_keyowner = "MTI" , key_keyname = "MGC-DVT-MTI" , key_method = "rsa"
`pragma protect key_block encoding = (enctype = "base64", line_length = 64, bytes = 128)
L+1gNguxvu6S9lsa3hsv3/w+vJ6YCSxDCPMZ4niZ9ZyaSau4cYuR3aFSffN4qZ50
R9QfxXIOGDwOwlDMU2vH6WJVsNQ/ZlcvPmxAEI2+zjZh10L0vqpt51rL3kVy2Bpd
/dJITD7zGQEZR+I3RP2wIhTshkqnDYTbbpvc3wFRav4=
`pragma protect data_block encoding = (enctype = "base64", line_length = 64, bytes = 11216)
oHQDbtJ4b2nrmsKcaqJXaLXA9m2tDfV2zGvHoFu3GxMb1V+MvjIFD/ghFMKMvFip
lewtwhFYy8mATZFQfZVITN8r0YhTzP7cZsABaBV4coqwefdfBOnLclBxjA0ao/ZW
byisn4ZHJjYkme8DLi/vq4Y+WzCr8wSmoamCNFh1zxZBpTs5m00ZzBKJ48KaQwqN
ZuXkIzfWjqaZN+giIoV2uhR/D1xE4LGj5bznUxP+QJ5X7IBW51gWK3w9BEtB+INQ
/kAMQdx83Lo39notLqSvYVhmSOk1XQa8pepgZt81eHoRg9nD9z/spREl6/ulF1Ox
aWSUuPA1ebkTalZpdVRGNU/rbzhgNl+R6g4hHYuwuk308IRbmy+SUyVjbzOz4dvQ
+fD/bfHFmVKmg7DZh2c4AOL/AdYhAi1qduFT/+fes2HX2l2g2JieuUivGex3u9pc
Njq06osypDDg05bfq41GVHCY9MaH8y4CWqHG+7gcK6VjWqNUxrVXcyAuYBlS847g
dscyQHRqNrwCQXJ8vmwTOb0RiDwOcse0iF8qHqgLlgoj9yxXvIVUh8sv2wPw6D9a
MFg3F8XEToPeY4kiRoJMf5g5K9YMlhzEHUEIXDHmEm8k6U/zstirZ0CcaEAU6OZb
iOBXzWnyvV7sbbNZLRM30E5bqg7KYyZkbpvUHirCJcLGZ2s4mHedXlkjqiEsSVW6
51XY9sqWtGV4ePTBpksWHAt5TwT1SdtXx8F2aKXpLfGyoEW2V4csknH7C/BoTJ/E
j71aLRUKFn6xlYcuWiEP/GQzpuNEoB4Q73tiRJ/lKepAmgBg6EzL3GubsTIQdZfv
w5vyo36tp4xef+qov7HAPUwf0urWNjvyAfeZfOuzkOQ1t2EGTaYhxWXkN+mwuB6k
PtD6qyboDqhxPRMPWuai4WUlYeLqRDyImoG6ZxRPmLFsdpKaRrJ5BtCQ2SNxUhxa
+WkN4ZzTEQDIcmD79xZVLdv+S2l/9t4kkMDpTMMkTrwlv3L4SIlIkGZAyZFb1fdg
wgef7enJqlBHWCOZzOb4+axeUIERPy7GcKxfNs7Nfum3hixv1F0TsjrlTDia4el5
OtIPVn7hPc4BhRdfV9ELMTKdoQCvOnNUH+KCHXY48M5foJIbuxLRy67kVtR2m0Xo
3y7znT+Q8FZCoIbtwHiPnbZp26dBoV75FgW9ZAZWJCn1LKR6pbjEsnM4U5N7sEcj
9keBuNd3URak+cHRmvSpAJYurKEGf25BX5Q8UBCFgpPh1CNkdzD3XrSC0vVLBNTr
axmOj63gfXEscLFItB7tccBX68ePBIfXJrvVwIiq+oN7wHMa/HSkHELiDL5/MG33
GXyfBkEwreACJSlAmjqPjinxqVxA37PBRwQ6hEbzivxTOuxt8FdrF735M9T/to1G
43V78R7pvjMynePGs/5ThqwPQnpknoR50NTM2NxU/fWgYulCf49cFwWYxLCGOGUQ
wQUuHv9Oky2weE1SHastQJ7RR3Z0p/mlRzBjA6Gp+xKjLHJZk+7d4uqGAN8INEwn
I3j4MOpWBthCwEsoiwmtGVG6IFN86apwIxbx/nOZgTFnD3DTec/hlJ3mbAV/ZCVC
0Xw3xuniGL2wSIF83ExAeJtu3ADEdL4kOKp/frFedlajCvLQOnOztCdGg6oLzQpX
ywon0pxvR/N41JAUlukzXMz2lMtJO4Olw+HPiDztAl8IbvNlJ1Q3qkV4srS3/9Lz
K3qOyRnwrSipLOTd9Aa/6SMVO+j5xcQwvNIS0ZE4HvZhPhUBQUszNVP8XcTxRI1y
JhO5NU3JhWa/CjQxLSjVdVztsSPEjOLkqQ7Pas8C7ilE1tIbjXEyaMxeIVVa731H
SHAmyFIXf3RbJ6fUgQejgwgDLC+C29qiYZyW4CBGMXn1w/+5BFcUSJbg+05NKaT5
W6BVPGmHaJt5fvzJ/HcMTCojdn9nskBuERSFITBhqcgysCrcLFOE3cNdOIU+vWBd
g0FRTNr68/hjPhvlAzxES+o5qfdhnWgayjhCxCP/y18M82y7ji9tZrnjoDDBMEhd
x6y74uJSS55vybu3xkmDT9g2kcTZgnVE97Q2eFSftO4PG/9CZnIrJjDhkztPyXZ2
k/DhzDpC7SpjR9kDV84zthJsrs1Pmou8FNlxEYyfHOEcYy5DBKUK2YPgjltqRCyY
Pf1VoreD1hh1Zitr/G9lXxAhJ80zOiS4bmryJUXIpsYiCzpLDz966mLE1Gx4LosA
CkhQZ9RbEjQcLKNOg/KFmXrwUNPRVm4Uh/Fhm6mguozzVRpwVFP2F5wYo9mjDEaN
HMkFw267DTh/PxmIqkgR5F/w2cdLp71Gu1fFzTK7tIbg9bosLRD0ApW+NqcixfKt
cmBwbUMmA6XztYUSY3AJkpgdvGgn+8MPUM7sfjT1jbdh9pAGifGgmYcT3mMjwgx5
bw2s+9f3JAkwComoYhXDk+KZIPOtfcjMch4NcEYBUjOWGLmFrYAmQa3+cfx1NlbE
9PfHUyEQTccSPaPl2u/Fim+HOM3z2iejM/epRzw02HMN08/kdnof0M1zMjyKWUYz
A+0weJuyvhYd/vVI4vTrdJYgqQWs//YvzjBArfFTmjMwKDcZyEIOuscC6KGCma/A
ZeibTFawBn3kFH2z9TlcEh+PF/nreKz+iYBVejZELqwD+7BOs26inptXu/Bw2F19
N+bbO5bO1eQ6BaFjg6+n2rMVmg9V+YigLxQ8sGKtYNzSm4EvIglUbcq3jJgIFXOM
2WX59QZi4O+IntiGHzFM835yZal2WfeElETWwNaNrryojyprxddVU8ykBke1ON8Z
VmQiW1ly7O8ikGIZioRrr0z+LBu/s++qWuka4njfmPY9qlYH+mtTRhfLKv/5UuL9
/ojOdfuWO6ARsC/3tN2q3KfhpmMGbkEVchWdNxRA/xjmuxOKdpFVu4WNaRY4fOEs
PCzEMIVX9mKMmwiGPytQIWYG8TjZ7IxCCjENEV+FvK5lbfYRewQP2IBLnoeeejrc
w4OvARbKD0IU4J05n/qGdsLeGNa5p5h6pb5VzxXpHqwuJNR0+d7VCJ3KWDxvH7h3
xwvrTi7njB1IOCumCuJdOxcax2cBLa+wqg7wsK83FQ6NVreoxX2/4CHlsARtiS9Y
mhT7w85llEO1oym0c+wVl7gg7SqJfN9vpHhOswY+X4D0N9CgRrzDaWDEPCDL4pug
0y7II7l1osMwmLpx8puurpj1Dj5wkNHHI1XFK8M+Fb5Z5Ug9ga9XrtQDZmdDJtrZ
P9B2aP6DzlWBLIaFuWSps8/RWcrXrRgBbkBwEF+OO51djkmaWzB0HTpdwlYJ2dJE
2gWR+6gxPeUZ0db+WCHEvR9LrlnYKZcFqK7PFbKvA76elRaDhoWdkJAzhLcz+5L3
QAffE/4DkmVggh/NhI9eiSJLNe+Xbti5uyKNYyfnjzOo9SxdzDPfSPwG9zbutNw1
X0x6qwu9E9vUN4UtxeNp0qG5s9TAw+XfFYWNEYwVSlmhblLvp5PQFLn9xlTdaHOi
S4M423Kw/sKNCqgQTiNhmexwparWlSqNUFkF6qgvNlb9Cp4c6xpIB60STGeYk4bp
R1U6bYniILHD7JaKdCmhArj6PnVARcDqxW8K9fCHn6VPfzY/ux5tYpqZMuXG09g/
ELkj5DjAdJb0BZCO0FkoTWvwcWvlc95kCamqAIfGh1DTaPXAxSoHXDaweBpeETx3
haTXVheIH3G3L+bqK7Vv7hFmd13ddkZipAqM+vhtvDXCexZJA9Du0K2gVPahEPJI
Y/FyARVyU91E+ov/tCIiRYKs7Q0KPy+rrm2aGWeaS0wRHcoQ0mjHQX5kPOi9ORHA
eQWedxA6bUEdC+kW1GWhgR2VBa/hwglZmY9RDykcIZHMmTHewZ0HT5F6tbP2EVuh
+rNa3wQpj3YUaEmeF3jgjRxmYHAeu3EpsM5BUF9D6AOBnga+PRBtKbKcVtYn1PuI
83yu7DXgrpXz7Whk6qwNWq6778XtWY6K8xuqBtdpEhrfHC0NWBrNvxIp6EAOjYus
PFXNNVYdQd2Mykcrx8W3eJaB3Qqhj3XUF9+n+qusshGR4OD/jV3aBCFNk3OZt9cx
FIbmFdY6m4jZjMmIUSYoRDIwuFRc+oWW0aAhGTkRU/Y3aKTo3tBr9NN8vSOcRZtO
oYnePqckzTmy7W7BLYDq460+0muhhGArTOrlmPO+ZBqDkJjU4UZuJngntrqI/neM
lCFIoYlaTDsAoEz44rrSFP8ZPraiytId7rq8dRlIxg4BzqnBcbvSPZC7klKE/I5L
mAzUH4+wGU2qspoI5TvoSNvWo9lZpI7nEb0MhIJtDPGzJkt6rP7KHkz63EbGo1T2
DgXaPn6pKXDOe7tfjOx9Sbo/4/o5soqgDv9vBPWVOVGu4V4zZekAFtQlhX6anddX
RYqycMBG+oQgjhswYektjAuRTJjAOq4zfh3ZbaZ4MdgIOA10tE/0Qu3cuEr8Lwc2
jYojks+jaBYc4MwdUq9Uw+5FT9WqYKa1NaKPmIlyg/5cLbOfTs/LGL7HBIW8oaDh
7uJkv2GobrTW3XZc/7umDWo4CJ4ndp7aCCNIawiVU4nRqRsZuhG35nG6FH07Kfbt
nES7MBC6jbz61MfBOV5BmoMvtkCMnZUZ6DfF6IwcCXMDWqjpW/8Tl9uYcZOGMBhu
XROc0QhQOR2ayr/WCds9fpDGLrJdEJ3aalbBgAAaklIcG/IGICz1NMssAuJsZyQu
Sw8kUw2P8ksa76Ys8P7LWb9Akp7Nl8tNqU9kBC59FNW9DWpbvdRsAHsLYQxDyWS2
5dCZcrprEmQ70Ey3OzbgjQnWL6UMHf+PSEgzuVTIhFn17r56JXDYxofszEsBPJsF
Z5nR2tMQ081zaRE9nJXwqTJ/Au89k9Tv+z8sMFhm8E0PgE/hc8n/5Xov71J6WP+y
kXW4bb2fXZdn7+nlW7uviUUPzAV/iqe33n3W1heiEqO6JcGBm8Z+gJRZRiznhYfO
R3HREGADaAg1NasekosaXEvomgxKbaH6L98nC4EqPaWU5o3KVcsrVwa+iEsvy9bC
f7RSQkNlkqKHrPiaP2dZdtqzZjfQ4eSWMb+k+QRzbou8Ug2taTnt6v0SIBHeTHnu
SBAfqhZMOQASSpdShjDwtBSa0eHl0QmhJFihJsy6pZwJ7pQLgQLxSchv0RfEhTHQ
xgJqKG6rGWTmZZsdGwVls1uiFa3ysQCHNHLrNheQ4xoj6JeDopZNLyxG04AS3eHn
55wctcF/dEPtW2xAPrYNO+L3xZuIke+zJ1rDmBly7VGsDmIIhWdN3O8q0+yvZHd9
Tuv4x3eJdz7fOAKbsKNCdmllxhn+KD2fs5ooHcd2Df7y6aWTdkUAVwDtGaPBgjE1
ML8TEv2W7m+KhH1fs1K50HjmwkS9nhpUlv1QDlpdZKv9f68MUuoZ6qyLCfXN4GlL
zEqXiCBKnUxwQruetxdCGz20Wpms8IFha9cEISyU23Kr4hvxsOtB3JHf0VZEo+Ak
Oz3kqeiEm/Ee47pOOmCa+RbEGQdHqgn95EBGJO+OmWPC93DPeccrcl97A8t18Vj/
pdc4wJ9Y7frWRHvFGqBhY1fCBvy1j1Iyq6OxZ0260Xhm/U+WVnonyRSO7pr0yevK
cSMBpOu03RRZnfP2D7vWlFClfBQg7LCAu0UIoXwlFm2v79+4mlBME9f3gtgRPPxF
ZwJup2lJve0hyP9NxGJxGrXMt2VLiBKj8gZOG4nPUiqwbYAXOrpQSj+x+cFbgKu1
LJ8hU7WQo6F+TFkl6QC9M9dMd9bXILjp2yWu9jcpdnFxG+Y+s6dSbJrdMf3gKRBl
PFSxMWdIHaAljyduakImBZ37oTIagpTaN7z64dENbxyxb116y91KmCLSne5Z9hO1
7ZFzriPva2b9o7VptpTE79lmNrBq8aGoN7VEaTrCOjUbbjlZeK9eLXctAsnQeON6
TbmoP5paKu5cXYnrwVo3jfdKDqSLZhAmpsBnKSEhjA2mN2CDebMdxTAOYBjwWG8s
vH2DwPjMiYpNtZ4CD2GIMB+zeK6LQUoIqXeV1VqZb+BndFyPzBMzLeMlHLW3riCe
bYo4ewPEfSWtw1tuNuxJA3O+0t99VhjLHQeKwiTcgAMUqzCxnA6WltDLTo118afb
Jy3uTQOU0iHhmFGEzviFBjAK2NtJGpBKvWR2B8fFbJm+VqZYzcNkIDCCIY0F7pda
pWMqb1ktvzcS2saEgwm4Hh1lp4ECP/xRdsA653KUha1Of25rTfyU06PSiO9ZnJP9
P6m14buVWPGU1x6CXfGnHm/j5hK0h6WqT9o5EuztmNiw+8d0gq2fBev7p0p0KywN
gGY0F8HZW47+FnqBfBmQ61ky+pTUYzSYCW+VFKnnJ3TESthTi1jevc0btPNpEIht
mxTrTuFqMrnRhdOjpiz7JHE94IbTUx27GSzIuddyNtdbohSX60IYqjRHRxQ0Xet7
OgopaxWw/hSyuMGuIO6GG70G2+fWwwiGaOTuSvSYvttndoXEk1LtD/v56wMrUwTO
dErYg48TGnCG85fKzVOTk9Cc67pVbisKkDhsqh79Z0OOXqjjcVAxw5twKZAa2BT4
OW9jeIoMFLuJPvQxaDwHZJNrbLLh4ZoyzeaI6YIONUsPqjLPLMUKFwoe5EtUkgjP
diSGLeviahDHZELpUETDI4EEjSXHT/76DGYfnttE7SU2mRCj7BnTzW07twoP+k8N
8Y1Rqe3bnTS7TC1Giu4IVStk+GZ2bHzQcr/FRVTQcQAjtNlUD/CcPrQE9vypQusE
j+7Pf9e7B7yL3mrzhnFuOGR/MUciwNlxIeWHGTO/n3nFL83MD3bNFEVrxDpBhmGq
U45Dz129B/Y99gUU2IC+bCM2sg4XEFjhbSXqTqshVMrQ6RCFUv+Iimn2JGnjD24r
815meljZlw9dJHwUks0ogtpocMHhbmzIUGBRP3//AkomEeVoTa6eTDqOdHzToQJU
vHfxrv+yq8kJCt3ktPvYgEn4F7cLFGrIlvj/37aYoSfSlVFrnatBz2i/pFBPbGxe
eEV44s070RheY9vUhPxNLgP0aGX8zjCKX6nAt8hGNlvKEY+uSWxaaRVReeZ1BQ7e
snWw2iyrjoMrboC1bAtzWyx+q/esY2DK55V2lgMWgFm6/oa+1kiE17MdRRwiiwrx
5Cub7u2HPrYovZomMmkqWIdR012i2kVDma5VY8SxLIRedeqHtnMwFatoNmokI9+R
E3WuCIFYwK/4CHlRKZHovuwKGvdLbSLvdut9qdY0JcUP7KY88sym4g4pRYBnVi8+
Nuoxmanf/3kcPjnNku+klAfC7mhKKTtg+z+MoO74/bdfM22+7g6JX5BX/s+kOiDL
e/vIeZQFnkOPzfoaymF0SoOGEuBzHMRE0752JNjNMvoUlkv7soHtr3PGJAUq4cUX
Hkn0sU0rsgFDalx7QcpySpUjJ/wOsiQB8P4QFkn3sKk6Vb5ndoq1y5zHLioPMFef
igW6QoGxR5r/SQovFPGSxgHG55rTixzXw/HjnlrMfFCoQz71tk4aK33NrfNGWMWU
qpgQZU+k4nGm42R3Re58HGHoUic34wgf4AD+Fz9GN+L6Nb23S2FRBrvG2Rul6kix
RMtM07u6awX1/b2hnaehXPCOcjQrQuNx7MMrfg/teq3ldWC/XmJMaQEJWdYvnsek
jyyoAu7aeecPZ7D2YlAYM9cgFpG1QeYT14vdn4zsxHmuQuskHCXaZlqt+adf9K/3
mAatgQ2BrJdAR3omnmUl8o6xoUit8gUOsA3IuoQHbpAKO3lEnI6Ttn7l/PAWOjVP
HeaTSrwDQ3nr+9oXqsVeEblX/RpA3AjAGtUN2L2/XxtIkjAiv7cJkzVm+OSmsvxu
dSBDSLBMAnRZ28kp40MrCWOBJXKQpqveREbeXgipfRtWyT6ouOw0/iNIJfxph5tQ
eH+G9jGoEm/YM1MoW3m0PGlPXf9ZOPzJEiLXJQbsbn2rTXpS6k8QSye6oQ4oJXf1
0oEoXAFuPXhuiyi73BcJXLlWzikdAzRK4NtdOIsw6MD3b2P6L0psp3qMkjZrP5s1
K4l0Wdp9xYDPaqFZILfrH2jjMk0h+FWEZeanILqmN4iykfx8PjysLIyWqdHWR5mD
+/tRcGbVHpx7+iy1J1hpHkgbsXuGdyyTGcVIWmTX3xe3CaZkwOteDFVtN+KKEz7s
95I4B8QvACf+gS4ATX1u4LltLEqu1PqkjiwBRI/w8eEuK4Jzt1xmNW5wpZYzNwx7
IaxmX1f449hdrWoZ6pTxC/otCcYFBhgjGiXRhLwh2EvZhlkwdEc/SN7TedvZOHgh
mYwxGZl/0YVUObv6Nf+02xYjtCSU1nWfuU4vnmVBz2QIz6QctW891gnUoEaOXSWZ
7Yp7Y8Oh+SHsVhQAVbepce/aLRNJhS98OEAZZu1febrOVS/ta2EUt5AgHFl15lwL
j3CraNPz+8+fB/p/1S1bWs9JiDp7fFfoWTS1l0iZ3YwJFlc7c02vsr+LQRYnvcW6
CBjsiO2tl6mHYzwvk/V9oAfx1z8vrHkrlB8vX8I892jCjEwd420mktch182m6Col
YB4Ez2jU85bYpJTnbEnfHjaDwuE5mTL92SS8YXHWNO1nq6Foj0OExS6Mw0iTW8cB
oz99okFW8xoqQsDglM1Pl8ZIITzkxSrx7u7OaPhNVAufLwN7RIbVZhOYXXLQRj3p
wSzQZrZb3ludk9ICNC1hDW/9vB/7TNbQYJbbJnFVoHg+sTJeEJ4IYpvI4qcjN5Iz
EP2SYM0dZPgMXeH32C79w7iHgevfbFY7nmTyr8iUmFlbzKMAkTW4PdesvQO2KHyy
h+Ifx0aBHdpnjziWp+wumua13Kv4KbgnSTPhEOIS9CztRjcQQ1PFiR859JRx3Os7
agFLbU5xMLTka46KnmoMx7JkVOf/+aHuD4kPaxcuo1qEYxhevcuQNm2MaTSBKNjf
YayYKx/8vwsPovYjErpQ51hZ5f8g5yX+Ks/iOBiEYNDaJRB2UZjKR/q73x0/XGae
be/gbrPkhdgwJvstyq7TzdNTKvceVFYlBWl8DNwA4BH2fR5B83I96WXQMErlPI++
U8FIiGGOdTo3T/xHbHIliTH9bvxMHwpyzhRMwbalMUBGBIQ3RYRSyW2LxXCpdyqG
nJcS+sHDO1QLvNW2wMSWBQq2wOYHiuQqja6DrT0CzXFZzwL/fpVVJ/1iOuJ45bVz
S4+2p8HZZrdrauz7GqFafDXp0yXrE37ySgk55CUg025k6Tw0uRlEsK7LblGY9/9b
+o0XnheoAEgJFjem1YKXOLL5t+FwuNb7LKE3d/M8uA5XfGkfGMrz4s67SRDN308G
CwpkDAjDR3AgwoL2CZqm6brVzhdinageT4bCEIh6SoHfROd6drw25MAIjY+1EVLR
rz6n1AgHDLmYIeD2y0pkeXbFNCalztCOAYQhQWnCtAvolaJNuRMulWY6JcMJfT8T
dVv0wjoeQmURRdotUq22jjjiGVMa6Xs44pVIYTuTA4xnPGVFVAJV1fpoLA30uBQf
attua/47eP0Hr9f4SqLpRTEsxjjBlwN0vVxcPn1G4ZUuhLfmepBLhaDpvp4/hCTr
YpBivM6HCbfs2MK3nd0mrojnhH7KbC8fOG4SyPYA7dlrlsoTQAPWGaYKmtuS5xql
zA/g/uQ14AlHno4nWpc6CMw3iCuFJ3iqOFFPMbj4dKW2nxeVFMZONn/kRIe8ujlN
KiznJav8dYGcDhXf3yUtvEuhOVlPDX/1Gwkyb7tnfRqJtM5cyKIFGQYDMo2aNREK
FKJrOiYc1wxNDXIB0gmx1dCiSzMjCIQpsbtiRDwFXjHrOtQRtuY3Q+kCS753ZbJ3
S39XYoPQaYqvttwFnkKpUrzRSUd4v5yWhaZHBHuhwDjvi8Cm9hYK2GG5fmsEZNdP
AKMoTXoIRP+fmPgSNaNctUA/hLTR3oCQWLX0g8UN2lAzRXUEa7psYPaMhm2hy0BE
CEdFTIbvrpvTsfyBfYUjkqUD8OhnAAzNhYgFPljdptMBu0Sw5Z5ltXGm63WFge9j
aj+CW/89izcliTxQ3Jhm0YAMzR2RDA9/jBSXC4ftlNpU/x3JisfBJZYWImiRj5G/
y8e7oeR+pNXO8fGwGAV7rSGeILUoq0a1DTEz/2JKtatw93103SXhMw+5Cq9ms723
90X6X3yZ7PaJQdND4ZwCpJenNXe+2Coi42diGLKQpV/njrMKQZi73wFwfT5CZuSX
YeBKVQClce1eXUK+7pDecT549GNDAJHWRKVThmy8guS6txvLIiJ/o7ofWxwkeQZ5
y46Jw5PRev6hfibXyHVRUYOm08zklfS6XAlOHa+B+tgUGYPJ+f68BykRFqWZVGQJ
hFbT8Rf2ThkykyXxsQp8vm0H3mMJwukgXPT/0kmSfj/njuK9oARFgIKNVggkUkRi
/dT6pBbZLYfanlmB2TvInH2bEef6zyFgdXx0S+B/RpGVOJa5/vKfcPMINi4u4gtx
oWNwYmgSQMNhq5NX0IdQcX/Hp/BgT8u8GRNQ5J9GKgrYuziRljkyGYqp0+CGmvDo
OCkHQdE/Mp6Mp85xmiMtZX2J5SaCEnidWvMlIoqeLfee2TX4xuO4hPsLZXAdYIfV
HBIvUzinI4UjuLbjHr/9pp3IE4vODhH25j/AYtSDVNSOBKhsQuOkHJgkOt1SOIk9
WX2kWweBsKSpcigHQJnzC3cMFf2ix2PaMor9VUtgtIpFiDIkmS5Wgjh5CGt9OBm5
Z08x5+3NX/vs3sNfRYfyLxofm8uash2CxYToubJdle5yDIF5gW2QhYw5sz85LaNv
c6LkKJLQ6s+cpVYjl7wdfuGlnBrnsoGJgLSBplewqhArHN9MO8EuuhNPA6oidqpL
ZC90/7Nnx02SYCFpwF4sm25iFOxw+MrI6jkSGRGeg+HN+EUAmc+5RXoai81oTXmS
KVEtKxpR/aZPFPKEhp4GoS/SJARU5Dx15BrYFIiYvBfNX/UhypWUf63aLzLJKqfW
XMrInXfuALvenRirrbef6plwuBTMKCPdqfh3h1vdn525A+v5ucccW9vHYbOKlUJz
PTCDH0I072KxacFkmCM2RF409V8wsoO2w8Rc4i9IHoQFGXhhFf5e9bxCapoCFmay
75b67wkaLghRyB/Y/cXLuUaxQ/f6GEHwY0+hSBJhyApY3R3QtAb9HpGVhxzrKof+
qqgoZFFuJRygS/XoF8WvI7/K3Du2AWFEIkcdBP6G/tpbyebTMdO4ag1v7p4x0Wzk
ZLYMFbhDLYUWZaLqto7NTja8PFAyR8Wbv0YFv1S2XMOH5UI3tGvfqEkdZMRVmq2o
2p0715ZYdoA+UBq+oexatFSjEndu4FAiIRWey28QUrBW0wFqZxu2TCy5nO8r2C4W
U5SxFdnchM0v5f+6AJg4oJASwhLnwFuAlIk3Kq/tTPdxfVlHG6gL+BLCHEwL2MRn
08oxo2d/R+SDnapbYPIaVSJNeoyz9I/CNmzr84+bFw8W7G4yjAxje9aeEMRsAgmX
KE1qPyFv2/96UWBQ7Xz5ao4Lb+OQS7cp22a0iN6fvLQ/RK1TBfM8C7kl/3RTMEn6
bLK+Jzgu9OInHn5IslPVCKJXpHoJwcZRt7et6wl0YSZJ3W0yz7EML/ALgW82UnN9
4IXAKiK20GXwkIkUjulsULscQ9rjJFeKmAcHm7wBpNHGo5txZzPybhRHdq4Y9txx
SrrJTyXsbSW/ZMD4XIBkRZ7823qyq2srE2ulZnNG8zvMtkQVL5ixsXBqE8uwUgC+
oFqvysokGvYnC5UrlOOHtf9se+bLziru9NnHFQ0X1KBH56qTLdECanUojwTEqeU9
ElFq8gZWNu2S10eES1JzWUXT28oMjdkdEEzPRLN/pzXeUv9uw5/SSfl4N8DfYtPb
5jWR2wbpN1M0n7QYV/EVj1ms9iQVsk5W8x1nOAAzYc57uVqIQUcxGZUGW/asDbPg
82FGkexxccK7GBEgJXVn+HuAn6sLPoOi2IpXYMIhWGI5lyuF6R1ijRkftskMl4Zy
wtOAmEwdMmRw8W1YIS18pxWCq2RbF1vNqcM6xOciwYZDBxnNLvRn+CEjrMgt6D7p
l1LazhLkJTn3A3mu8VpleTODGlHXu8xGS4WdALOmy1lgK5zwVCW5X5oGNGnhC/3o
vLX6hViJXha5HddmdmdSmouSNaJa/eHMSIE3/elTU+GBGdaw38iMg1Fm9CepFcYj
q38ZFtMipM+QkjgJrrB1vRsjEfymyxEfZAQ573MCNHO6VL2J09pJMP/RU1bzRw3i
beMUTMV6vpVpNEaTS9JJ0YC6Pm5xSyLY7z7EropWsZatYUDUP+XfeWlRVlZw1YvU
/vaO+nFNHnmbO/wpXRsXx/3K2MQfLn4+RidXduaKcjbS9gfs+d0hBcQY5GH+GFPz
NSSUJ5hWOM0sBqGwjiqNLPB+qDwfXxVsgbU1qeIYPCUlalfCmrgKyrMy7DnOVVCp
eHtQfwb+Yw6XAq3VhN2arF4IlD7yUvKaiUU+BvtrN+pUG3XjQkCmdkwAifxnzx2n
t9ECm5uZ7bArxi4mB51dICOHvMWUDwtApRuHICxzshZlLs+zlfkcFpDYcJ41zATo
+jDcqYGgLYr6Q2cG4LQkG0hZ4JoaBQw6t8bM+Hb77UwmBVCAFajJLPY6Wu4mo72u
naaZLqZi7sbgmx6PSKtm3PRhyIAeleESpfbwcB+mFKHw86IQRuwbL5IAQwxgCE9l
25/8KpV/A7J1Gx0liY0umWxWH/FYMQeIUj83OfeNL33TQ6uJL+mLqXAXxC0e2Z3g
nwwHmPySLmaHa0B7GxaX50ywJSaN6SM3qB8n6G/0tjj7A18SfxqUOuuuEy9TO4EP
vByev0llvbpMfQSaNozbB0W4kYNzYmr7QJD2oTxunMCaTuZpMCFNC4kfi/YPxYJu
c5kDSmj4/QsPtcUeSSIkl753Q0exiCrCHyPWQa37GmSASArTZpcFVEAqFqY3/6JX
J32GIywM94g8IWmWMn0BegW4NduSOSsPnH03NpeC+uKdz5FPA36wTcE2yRvKl31W
sMHRefVq0XoqUYg45lCRPwC1Qhqz1W9cLGIe9nk/29eC6qVnqsQ+e0WHJMMB4Nto
3fAeDOXYcqiYLkjwrfssTZNT+addNDsxJ138pdAtRC9Q/OAioH2fUdG49g4wAoAb
rQvO38jV89BPka4baR/79dVECWS2BW7t+RZ+424gDFm2jLTcw0aexvloW7MjWFDe
MBRLi32GP06bgHWj808LY1sVblS1+m7IiNv39YSRspJu5J1BQGfIqwEufcsDt02R
b/S+JbCfVXg0rZ/8h+udbPYuDEFUHZNcsOHz3Q74wWx26IfVvE5LRp04krIoYoIm
7rAGXYZof4VqZGuiGosXPjiC/rz2SGSUKZ1rhIz4/Cb+pIiQ8de6ZYT/P0y4OgOI
DyJ5Nxqaj4a8QL695C2z+zdBzKFeg6gcpJxpVm3Blv0+LI2hyeV6z0E0KfJ0tGK5
RmMb6MfH9iGZdxuDWa2hglRr8uod1XJImy9rmdLhNmOyt93O5eLqAKUWOFmwDWkd
cgjlITeKxj8QeNl5R4bQhhsxZr5LrMLPixWqa0uFxsCBs7nyvPsBeYHDEtaFvFo3
2n6qzBQvkUj13L1nfT7Vj6F4nH103h6adVR6tvtzyXpbVt7GSOzKJELAeWnWuP8z
FQVsq0N+teH/6NtnOl+56w+xholNJ1B7dBWohELiiKdQN0YzlMjcYlBOGgibUfS/
zknZqBLMSX3EbnfFaru9YI5L8nxit+V32vqO9SovwmXfE4AZI471Ru79u71boLVj
AW9XqanNFY5MBMYeFeL9SWDwLOQGwXSw1avc2ELe/A16+uCYPqK7tqCoaxiqlg28
3TTtkJIQX4RwwnkUILwMoP5t5xLdVcMCmAIWrFsbWTlO8WfIw8IEGbm68QoJ1UfV
zsUsMpMst+uCHhwBRb1rWi+GbgWilHWw9pzuo2oH5wu8boyotarUQkp5iw6MiGgv
wIvqfnHMKbC6HXwf5IUK5qEOeRZ9rnm8b1qMVV8F1v56SLi/rRXXox/OE1Q2HnzN
z/M9yIHYS07DlOcwoUSgQPd4eTC/1hw1rRMe/TC7egwcRu3XtUrn2o98bRRpS5Hj
ZGDsfqkMdTpV7rKcKwR/btS7f6lfW6b3xQqtCeV23q91/gZuwE4TTJFrMcMuYgx5
SeHRdkk1M0SvAjIsQIiFcy9hoQhvYM9/YRlfJ9db12xSTfiL56ibi0Wa76/4sq1n
/leIOQv/zNcEnPYijWTwUrCPCdNVnfwuiHnG32uBQd7q+M4ndOTzNmO0PdicX/NV
/VjBfJPPPZXIvKFoMWaXBDntQCIOMdlXu3CE2oPn/zVOFh4xVpyVsSZNrW1LOTRv
7B0dwJ8w7/qz6X/+ruvkP7yObUYdxPDwyLeiIvOZ02xWNWhpoWgXZ/UKaa9410tS
Khu7Z9k5PF1T/sH+w5pc1c+xqYWmFnzSEdJkoobTAIZm6l9nvmtI9vGWkamjOTwm
W4sycx0EzbdkVK7Ba7nRk5y1grPE8sqLqLW6+P3nXqJ9d5xGhdyk6y9oYCOIdhx8
Y/mHrvCCG6RATzODC3PMcYzjyBolFGwEDh0iyVPklTmw1pJyA3AHjbq/BwLxuNXO
BezIPulOwLGNl72xta1R0oxEm4W6kHQVgQOnoWMnPyRli5otLfBqOH8pAp+X2Gkd
MYRvYreDgkZrlkMdsbT8ZuMpC5uSw+BKbwUcnvKQEuKloVJYJda+9R0vXX2RAD5/
xM2yyr/zxl97m1lxyFmKTop/3CFPZ+CHVIgxzi2SHj8wcfs7EuNDbsBSIXXGj/Do
c3n6TeH3Io1WoDVwGNR0ygh9JbVvIeM5MKPY2pRm/X0jlMssgXrFcMLj8Am4zybk
D+T7SbNZ5gR4UAPYurFomO5HLG1YwKYcj+cZGYINIDY=
`pragma protect end_protected
