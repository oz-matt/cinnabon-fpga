��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o�X���3�k���(cvv�����ܤ�5�֖���\��i�L�2�sq�fD�� �wY�J��l�̇��+�WZ�<�
�m���XI����.6�Ii����7a�!BY�r��XR �{]�����A����-�\�kѻgOtt������R&T��[��@I�3;:�S�#\_�F�2z.V�3����N�(�J���%y-�ͯ��Xg6Q��.K/�U��JJ�_�Ж�5=�����:n��b�>'�D�H'��M%ƍJf�~ �o�oTasA���	}H�+J�(�	�����(5�q>ԗ�	�q��������R���&5�-X�#�32Xe�"�L�z��.R�_(� _�G�u:����I_T� ��	�����-.CC�<�CW�q(��6�ڠ������`Z��j��x���_;�hZ�(����,��,�=#�T���v�1�CdAԶXl��&�v�>������K����όR��9�0Th�L���Æ�2%��Q�s3��Z`G��*���� ���a��:k<g�gq�Crm�$T�U[���x������+�G����.���-9��cM���-Rka��k=���7Y��.���I5�w�/��6W�읳�1vS��[i����m3�:�tp��R��� �,��Bf�4�&Z�ը��S~��]n�m�9ѝ[m�-����:���YiB�LE|�3�eW<��L#n��)�Ҝ$����4���4F�~�(�������{f]ǈ$h�v�X㘅�.�����X��%)�ah�"������z?cP`��A��}�~�6��Ӑ?�+��_��c���3��FƤ:)6��f��>Z7%]Y�z��� �.+d 
�$��|�C=��$�C+qo�(HHq�T��~eЩ�hbI<�i}&e��1lq���=��_+D�>�W϶��X�k-�(Ҟ� v��(f���U
u){e�Akb�6w۾�(2��-��whQc���atx��0__~�vQvg<'���ܨb�ch����JaG�N�,4鐽#��x!waJ[��(�z�3L=L�U����d�:���S��f����u��_X��m��[HK(�U#��h뮂�3[�vW_�Vh_O�j�����1��vW%�>�X�!��o����5yc���TR��������k9 �h(���T�xRΪ��\$����E���yR���:��k|*j�9�sd�?���a�n�k��x��hS3\�#�86��v���ܚ���J��vd�N��$Q�A��1D�T3U�S�T2����6�<�����v<cDbn�,�A����~
��d2�-�t�������;��z7�f��� ��JU���:�}�wPj���f�>to�81ss���S�]b86�6��� %ԝb���ʐ��?��������:`(�5
�u�h8-0�����6�W^���7�Ys��~g/�*�8n_H�7O��e��T�\��A���`er#����9
jEK�:�k��淂��aҹ�5�M׸���C�!����G���]�$ ��Y����4���h��=���	�/��{t��}�q�j�e��D�y!Rq�2�y���hF�\�����c&�H::�}W5T2�7
�s��Fl����Z��l6?�n����t��e��f�@�=��p���t��l�u��`�F�ʜ �($mg��xԩ��]���?��hU���|6-����gy�s��#�9ً�eɱ��AN���n�%4{*���J�5��f}��Xi$6U�a�H��$�5�eQ���"�%�ʙ�fm�GT~�>�|e������ш�.�G�&8x
�>E�K5I[pN%٫���O�
\���k0�N���YC��V[Vy�/�{�j�/"?<r�Q�O�3���c{ ���Z0���+�N��������G���iJke?�A�����'��@n�G�y��s�q%�$�,v;7�0[�O�j�����dd�@៩��U��$�0�uSF���P��$�U�/:~22%�8MP
��\�Hg$�M��
��x�򶩹�g�n8\�f�ރmv���Kz��Yp;��-ϱ�Z�ST���w�-����&�ު����0�s�Z�;�tx��nC���{�j{v~�_i�T4bǭ5��P��v�o�e��L���tMY0=9����������� �h���~:sh=a޵z(�?P�Y@z��=t�g��)�Vъ��y���,Ü峆����1c�ta�0��e���YW�W%���/���M�(9"�+�z�ƒ4�&U�$�.��@�Z����5B9맶�Ǻ�pē�5�?慺��.�x�F�iHm�:�ɴY⡻D/�E��Os��b�2qZ�~S�#j����v}�Q�P�D���(D@��%�~�P��;u.����[�7�2��"X�"�}b[�K�0��5<-C�&�N����1sc��(���m�B+e�Z��߷�����-I50M�<;Q�{e�.����gq�z�Z���5�	��	�*�����O�i�2	�=���M��.�ǔ��jJ8]�(!B�|T}���B�(!�u���Rc�j��M��.�*����G�3~�������aB�F�T[����tV������퇀-�h@�E%��3�]��nvc�� ���t�)
��v[���ѿu!oE�F?[fJ��vq�L��K߇�(�w"}i�)��`7AnY R�灴�S���ƥߒV6���^Ű�H�t��x!�j�u��ߡ��2%��&��� �B���������u���mbe���U�Ǩ�S�?I2-�|�=9����*�:�@C4t\��K��է��v�iÝ�GV��'���$���(f�A�;]���P��4���a�`��[�%�	}Ql���?����˅�;ONM�`aH��P��52p$��*8�	,l2>#ƪ�W�@��e�9:�� �W�N� �H;�J�*��=�jn��X�J96GjU)��?1x�r`.J�#Qƨ��3�1;�ʁ��g 4�l k�)�Y�>x3���󰝡�*|�ό&s�2�{O��VT���j��	C�v��D��?��Fh�Mp+���Q=��ׁ�69'��
f��v�q���r��
�ޭx���]��]&��eZ��A�o*��%Pi��Ȝ�)��V�6��,�-�Y����ԄA���� :�▊+p����W;���gN!�-�+ �j�/��
�1H-�|�0\��r�G�1�.>�~��*'� (�v��HW̭5$�'4����̛ih�gy�Ǯ��ci��&u�y���!걇���9���E� �/o��dY�4a!�|�G�l�� �זX �^=	�ʀ>tp�9�To��}�dP�4���J�P��:Y��4qzҞF��T��|{�%�N�C+~sDh�: -�(�?�tsk�q�c8��3#��S��{RG�q`��Т�Ig�<����t�r�Q ���ǵ@8s��0G���ъ$_�3��L>�v���׏�}����f���)R�a�pvcg��nŮ��+hQU��a�zt�K��&�9��4��O�`}���S�W�=������r�Ql��A3���P�7�J���1k�BFn|��%p\W8%��T!h�1$���rJ>ȍ��ߨ(m���sr	���M�Y�B�q�ҭy�L������� �B�Lxy�B4���{�?��鄙.�҅p�+S�`Fcl=J����'�L��̦��Ʋ2
�Bі�*���c��3�^��Λ_{}/���~@k{�WU�Y�v7Up�w�b;��P���B߅wr����f	�n�<�3r�$<ٍ�v�=��JԬd���:q���?x�h����sS��@�}���w���.��6�O�Zi(*�N�KC�Ռp�b�WCm��D�7ϗ)��^8v��DaLapw�oݣ�wZ������L˵��\W}�x~�*9Dc�U����YA�w�|�z|�Kv�&�i
��>�%���X�1���4
>��B
=���j[Nlƶ_�*M�dNO����� c��y��Jn�>߃���@n���,Rm�
�T���!�J<̓���j(;���:���3�I�w�d�7��^�2�l�6�>s�kZ��Y>�L�ٚ貸}4�c�cZ�c���搒v��gʋt+7��N�l�4�F�����r���U+�����_U���|�\�ͼ� p/w����^�g�M�'̜P&�29mg_2K:NJ:@U}y|�]�\���:��B�7��:;���Y>�dI���>p�(��i��D��X�ڑ$�}Q'�T�ŁNp������j�����f&Cu�%���Qs��m_:�f�՘��(���b^�$̑�n>�W���2?$ɺ�}�؀��	&�y9dik!|_h�S�;5�D$n^��J����O�)2��J��̊q��,t��֣�"���#�k_�ь+%hH̳�8��GM���N4x����96)�?m!dS�a`���qG���y��ۼ����y�@�2Ń���-�q]_J׏��ǃ�;�j+m^�='�ɭ�p� b�n����H�'�@B���⁝��o�t�|�^�{�&LJ^>Mo�g�g�A_�L�R�Ⱦ��ͭ1���T�3}_����|���W��.�}BW+�-;	n<{���lAB�����m͂nXG=k!�1C/�A���
�oD@0����D���L�Z�׫u��~bK�� B�����)&Ý�f��v(+���3��ui2��>bG�3�0��݆��Za�KU��+�_\�kX4�W'ڶ'8��)4���
yG�6<��:z�kD1G�ӺJ��)��J!� ���G��e�q�p�yA��i����(8B_��ap	Z�3?j��!���E�%��*���n�d������5/n�a��I��;�g�_�V�7�j��h���N��2X��%�,b�]���[��Y�
�̎)ŀ�8Թ�8�?�\������Eل��c�H��٥�I/B������8E�<���o���}d�����ݠ�k�W7(w�=L3�Uq�_o�G���	|\��[�1$�I����H�5Az INƮ��s���r{�4�fE��j%�o�ODr�ˆ�YR��� �e�K�D{���39��_,Ig�;P�+���į]�~n͞jgS4t�g��tNr�� �O���o2; �r��䗂C$17��F��.{XAp��WK���0���a|�D��	4@��@�n�!X�0ד_[xf����×����?�t����v6�9!y����j�
��&>v�(�+�P�ԹQU7W�
�ώ�a�$���[6�m�0y�8^�޻�}�D����h�����=�}E��M��{�['}Ays����� �e��"(��RX֦�	�{$�SJU?���(^���^'^H^��P�Ƶ�m,�ܮqGb��6���@CQ��MQe
�nq���+�o!�������R�����@�x1ة���~�;,Ϣ-��gc���	�q=�ח��5�ĲX���9]�'�z>ī�33A���\�p����c�u��+�dojh�1�c1�>$8a]��.�#vc�h��1��W�~!����|l�W�F0|�Oz4��py�h��<���2$���R0$>��S��ѕ�e;�G)P�]�;�rP2��9+,�qj��\T8�6�phZ����İw]/w�=�觻ymj�HT�Ĳ>�[��8p�G0���Q�|_��Ħ_��������-/،�h�uh��ȎzS���؁��X^�?�7���o�|�H"ct�A2;�s.d+�����p)�c�ݎ�a<�I%L�O!������E �u������=�߂�ȄܧX�=��)-q�.|@))C9�!%��PH2:H�R����|�5)�0�Y��?�/5Jװ[��Hq�����ǞgCZ��ʃ|Dy\<@�U�- �&}m\F-jd���k\��>��3c���ta��m)D(��&)5Wu/�M�<5Z��~�J݂�­�6�i*�G�%��R2�l�V.��ijA87��a\�ر�!V��1��-P)� �-hZK�?���D�	Y��H<��괁�l����'�2ޑ'1{��;��	M�uҋ������$�n�/a;�{TB�`� �Ae�L`G������V�'7�C�E�~\2��$����,��.�n�9Tj[�PZ (�L�0RU�\�t#�3�VFxg�r���0�M�z���_��Mg#��U�]c5��`,��_ʲo�KQ���)]�!-j� ��+͋�d��p���	�j�n�+:>�/����(J�ۦ�D����܁�t��w�';���]�zƴ�r�ۅ@9���͹}�o����(��)
��"��@�.5#�	��!�p	�^��{T��-r�PAj���� ;� ����8�g[��V���mO�2e֭�w&����R�☂*�]}��K��k{��������5fxVi�.�{���5��>�u`��#����?��*���B�Й�z��DDNä�'��~�@5*�Yw�w[�@hߝ�x�)��b���m_'�i���B��(��v��
�r���$�L�@�nע!G��o��VP�)�87��ZU����D!܂��aN8���y>��K�u��{��>`=
����]�3��Ct�u�7a>۠��Ŷ�0	�ކ	�*������p��Rli�A�Ep��R�ީ���d�"p�����v?'A!�2���H�p<3���R�av����JА��.m}��>fmj���]��/��'-kV=��+�|!+�%��eoZg�I���s��Ji�4��!�%��X+�Vw��-S�Ӄ;ՌqXS���3jb%ק�^iA��Ti�˸-&~�+��;A:*��|2��ru�t�|Cr8���浛�۫$	��Ԓ�R�C���d�y)��H��!W9S������wr��T�"2�T���_�s�C���d��zh�$��*q�p �{Ǽ�DuzQ:v)~.f���G�l�]}�E�u|�^�0�jL�Z_�@ו���!i�z'�à~�V+��&u]��<>ՅDq��Dv}���tZF��0� V&�48S_=	PU4I/Y[tl�q��g���*>�_�2�(u�����L��_��`ђ�8:>���y��_���2��eˍf��Cv�P�)E�:��ӣ�*#����'bN�W"P�j��>[ۧ��\m�;���6�T����[X~�6�H���)�72hI�aa-B����L��ݡ C��{'��'UlmTR&�^ ;Z\���eLq"*�4�Lr�o |��E=���8��P�%oMW%͑��F�_�LɅ���7\��n���o:�3:�Ŕ��^!�6��ƍ�������)��XyqI-�'����H�B^Y�F=t@M�;7i^�Η�#� O"���Wp�?ek��*|5�~�M6G�r�C}�����q�&��O����\*�
|�݄�هQ93!]	�$VR�- ��F�l!	�݁�z�*����)��M�^�|�rs����@.P=0����r��Z�\�p��vA]�$�z�KZNd��F=J��@M� '��G�`��j�)�C����v���V�nE`���8JM�B��-� ��W�%��r��34%�O:���z��bR��{�D�25���F3���]罓���Ne��Jo�q�Q|�c��pݞ�����	=J�F�����yp��06@���}+�c�d.�樃�`�Q�L�d������{�鄄���מ����w1�R~�,����x�~9�FN\�qk�,ʩV5\2��Um�a��8+z���pA��*������duW+w�IШkX+O󉲅��{�;�䐴$K������� *���	3���P�ri]�y�?���p�v[�+�(Z��W�6��n���S.�����/��d������5��e�e�Uc�?��*?�D��fbI�q+�ق�f�h�Q64�j�TI4y}��������ۄ"x;Ss0��n���A2�lY)�9G�ȝ�d}�G����]| b��[4͜wHCzqIaR�y�s(u�7�U�*T` �F��\"�ù��ZJ�xQ�	������<����E���ǁ/\Ĵ}��T����=��}E)O��y�����Y�T����c�%0��Y�R����&��Ÿe��\��G�0�%I���4(U.��7���;*Lg.�y;	sy��^t�����p������d�2�z�n�J�I�Qj�}���2�(��IF� �j!�kac����d��]&�Lx�)�����{����!w�Iɔ�^�@���0��ݛ��kC*�Z, ���ݦ�*�ߜ<��6���5�0�d�%{�I��i����y}j!>�yY��L\$3*�S4�k(�Oe��jI�>z<p0E3�[J�V��U��	|�n���+��¡)��Z��sF ��xKNm��;<�My8{�A�Z��_���6���4r?�2Or�P?�R��~
T�������aĳ4c�9�sO�s�na��W�%�'��( ��-@0�~�9N���E��pv��n{�׌���!�z��N��5��*����ҰI��Y2/�9Q�Wz�����)��W�Yw�f\]��?�ت�y�ry�(�,x�R�!M�{��;xA.a�	�z�ءGYp`\�	���֪YL'�
�{���=���i����I��1�q����:5��/��oT�]E�&T���-+y�9;ŝ���'.�F+7g�&�BP�����Pd��i�c�T�W9���b�P�4�<���߹Q.��Bh��S�+�N�"�+t��90Q�^B��%�G�KBr���6 ��r�p� ��c���S3y�c��\D.�T�����)�ɘ���y�s8��(ֶp�6E�߁��.�9���c��ji���>�o�ca%*b�<���WPt�Z�(���`���l�v㈿���2�A�á�	J�o�;��ǡ�Y%Y����2]�㫂a����!TmI���|KD���0��lsw:3�L�"擩�l��8���xm ����n�R{&�EG����9@0+��ez