-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
bjrWiJiwAXEkXQFYvPhXjikIs7RHMRVur4N/RAyoXP8t5tMxMFRGOADNYfilX/2qZuU8GOvXSH4O
evmz6dgF1mS8lrciFqwmssdIhu3Tsg/vez7Z/NZ2GwbO/MP6NLUor8qiUpgnn3rZlpZRB921QdVt
6wvLthAgsD3PKRfrCkBhAxpglGGYVu2F7fIfNrprKoEWxHgPgp/md1+a/nVKb/Ilo94ZFeNvg5NM
3kr/lMVSf4/3LZXQP24hTOk/mha+96ELtm7cfVWp54802FonGSXWSECHicaV8eJBxvJQyGiA8rnC
l1ZgYwjI5tLRFGgU6eh6calbI+XGTbuum6qHYA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 4832)
`protect data_block
M79ZLtIA/slhtS/gjufjbhN9bapeBwKuiFY8mNlH6xbEyD2JLzWH0JelJW+HHiph3iw6/u04ZG4w
aLFFA8Xbi39ASOykJU/pAnn3GOlywPRfxJ7gSjy9Sg+4jWjDq1JfxHIEeFZx49CkjWvmmVmMYfiQ
rTozOU6DbDqkL6Ub+j1chpxjs/q2MtD/0rFSl99zS9EkJEflEosomY/zx0shN8PbAeF4OAnnaBtO
yJDJz9SNgSVQ7lrm0tW1ZSAflXmUG8mUVw8Kr89t931EpdUA7yp4LeOatE1fjxPV1hZSc8ZP0xPz
8pf3My6Y5umLf5rDl/GZaUI2LDnLj46Hij28b8iLg79vOfMAsq7MgAiUMavhaRXz4kAMBLGVtQqH
dEUU+TTAYUGOH3se2Zeyn9n6+2dRAXAQPnarrcm75gzjHEhi/p12lV3+Ky7WHoS6JLW253l6323b
fVkpO8cdDJz7esvwV20hb873nF5T/3vaRuMCpLjnzjncDQAcf7YmkbM/g2rx5zxX4mZfDFISfO6f
0wDFAc2w5JaLPe9B43+hqIraDMkoUwym1PXST34fZNMW4y2LxO+X/wj90sDhUPc0jZ1UQ2mlRJ6c
8JGyddosD7sdLeb9tcHg5BB+WLAjPeVenHrLhUffb0wVOY6BbUtMkJORFIlc2N0j9VIAyFM8litc
pnmxaYpVsrKMi5/Xq/d5dgJiMLRb/fMlRHURouq7yHF/r1O1K3UU+plk9t+9P/OHOk9Km8fgmAfD
6q/E2nlFpqpb//hsuoPz4r4arFgK88LrGlviv+Bnkj+G0b3b1hBTu1Z3dMyANp42ikeZt+ekCHKg
XjcK6K1BGgIIHDTzsGbaZrYq3DEurOdu4jN8WYj6GAJ1me2syN9FRTKhqIvXQw//hfHFSpkpaz+m
PdCdfiGZ/9OmRFLia5WZgfyb+BJh9ABeyn/TMub17wKrhS7+CbYQc80YOpscc2KIIqaKiHL9H7hp
RIVza/G1DymPgAUO+HTlt215UEK+0OZ/drsHYJRFQXT61yKeReVaCxlpOSUUHSMczV1U+HxS7WY2
azezQ9rEexdJcxDKiRy+gIhql2xB9eAQSS50jNyo05i5C0DnXrjOLVJQYNPoWKbgAPeDslDXpbma
vonyxgqEjrbpHSFX+HFzqzkCJziL3aFbITHWUiAHOqGtyVZgZ3og122Jk9dOuuYI684zriwvEoTH
mPkbsTTFn54NmMUJd4wYQBotO/tSlkegE0+7YvphiRT3OWXXxCLckUL7D6xNJnD49D/hS9XjPQeo
VBji42pB/Ms447NIPaUsOjwNkd8RDuaS3AzJQMk1llW9uA38BX7Jpg3+ZbqahkoWFvrh+Vzm0EYU
LA1AsWSULNX6/MFK39hirrlyradfST6P/cbp7aTLvCeWeWrfM87C46PaTVdvGH9ihu3tnvNPEJvc
GcJHsJVHm8nFLuDiceTNt0vd2SxtKgcg0RGSIBq2ehB1/fdh9TiDDQURsdHhP1DUwcBKB/oeOSmZ
iSnMO3vgy21kM0wbn7HsHzGMprc+KecJOjarIIZTi9HeLHChm9L8JIy68onBO2lVNS/DiowoqMYZ
w9iHdveaxCUSvfTHcw5gHl8l3Rg7Ix/g1ikZyJs0YXu0WrGfAm/E1uwXVaGXotttyXZMhRyGskpo
iNq7AeXSRYAlFtdwgwBnR/4Fj1Der9Thav72d57hMU4zmyftEDCWpXhB7QiVJ9nkOD6zZ5q7Gs2k
cXV2JHx8plshS6/5OMNvgYwXuiMiFVzu5NrU+qf58FFmqQa06ipNfGi+9G14ZtnCb+sUKxo0nke3
agQ8C/rO7juI8Si3mw5vdlsvSyliwa5soeGTZp4Edm5spblkY6MZ1jH7o9ZSk+tJ0IXYgk496KDU
y2CiMEbc0RttFJjwjFMf5/gFU4q8dn+tw9td5nDIsgUP6H3e0QK5BISLXvHNvo2FAnJpwIEryCy0
5IbIL1RBrdoKaY7Dc1mN0LQ78poJTOeXsN6j0DQ0X/hgaGVZB9RSxtFDIAqNKVeg+/zI2HHW8M4X
eWUrISCSQIXn8tzA31Z81FpQH4Ihdk14d+oZIc9hHXvTnuxujUSBeEhf2Pi+L/+4d/KatTgidHvD
jjd9knarbdMZwlxWoQlDdBDAiEkMvQ0qLF7GATrIyXeLxpjDXwIvj9fQwjwRJfMxV6IyOEnB3ocm
JYkIhNX0qy2LOSla3PhMycpkC+MeQrr/br01tBgdRlPSJdjkfn9FhXVgwlrKeRELoNj/Zeoqs/qT
3AnSSR2QxWeIRqUwYcmA9gY/WAgVEMX9D3j8BXtbWJcWkdSzmhAS5vKOr32PaNOcOwIolNHP/ta/
8q50KGuzEW3e1lkum3q9lywQ1xcFr6NTfLzCZhuhXITpBE5hgIsD6cvj8apFzpUg2bHDxc865kLO
68p1ITBAjwP4jhM3s+I0DcPVs1k8bosoh2pdmwRYgsOipCC6cDmHKUGHEo5wLOJejGbwHzL6G5Q0
96BOaCxwzHAwtSyDlEBz5FK/dLhkcFZtMfLkMZS8hiO06CdIJbfrNzE0b7kKALkAhqMy0zMFzPuH
mS7JTSNvHYZOSz0eMwuLv8xOMzp/K/2A88AaGdrm4iMtjpiZdCsVgftgNwQNT2BCUOMfpMH2+eqG
hsvvRsg23+7NFndpRf8BVXp/ZFdU+NiyHh9Jx0ukgfa7MjtdaOKl1NlkhurN8V+4uO12B1/aqA99
vIzItA0KWM2Rns5zh8YDvHF/qi0ktCtZ1P5SQGpPhF7Ak0ZhXAE5Pk0lcO6ScEAdketMmZ6erEeM
+8hz9o9LCKs79BC5Qkz4cKD0atG0s/eeILURWdNrn6Nrh+zqKm7hbuOhSmSAAkXuT6M5CStSSBAE
USoMKoh81VbcWbuKZIPImoG1GrygPP7tbmRaieCyrPFYz1TmSQQ2hSDOU9YozVkJktIQ7Aod4M+s
KcUmmQGfL2UCTXSnkypvd6rRg/VMhvTUqfWjSfToSanROSThsRSshvbt/bPvCgsv653z1Mz8JwmV
1EtsBiSajBqT1oT4Tpz5fhHW3bjZOfDeHs3SCoZ3c5Ll6axzmVlabGL8Mb9eAW+2fNc7QZgi457D
56fiVOK0VfSIk7z7YYJSyQMu8CPi13Gdl36buQ5KNFfYJNVJztFXEj9NpZFAxS3v+zQpEG2Ufkjh
LRWyC6ngrQj7MBaGDoHNHWuIjqaj4n4AfHv4Xz4N/Jq13Fz1aNt6QuiZmzTaCjXvUso1ysbe4myq
yIRWBOg9nUIepTjLhAxx+7hfZZlVmH4vBWjQXfWrjiotYbUdyVdHJL/Fy1h7TG5eehquqjVzHmiH
1wJrQ0K6MHxDS+Bw6sINJwW+EEXQwkEdKW+fnaAmDjOZlLNS7WGHDNJ2B7ztfLrNuhp9n7KN3DhA
OTMJ+7Ta2V1P2u6lLc7jTrKeu4vWp7cF4HgpK/t7khUEmEIuRE2eqx4K3QD0x0h3NgyIvzLgg/Jr
f8muD1S5oJHldmyZZOiHn84R6VKMfyxv/nUDdr1K4dSBI5YKfTjoPqPG+ahJRaRUplPFFe1sSBz4
TYWO4QpiDOpkjY7vrQ1+osHKxJpcRmFXjWgAwCqEXoWqabU4DQ/61Pisfib962uL/au0JIwbDsie
7vSxboxv/7IV3Yx4FLlrevxeyzfbLHb5bVo4TeAMEe071M456n4/pHfCyNY38PisUAayUPpL45m1
aghZqYZq+LfvUrbJlZFRoa1fH23c34RxAtHyBPVGKHiVyxohDAjVBCrlOtU//R8bsTY9BhAvQWR9
6G/V9JELyzxf5CtE9AIfL+uiIpMwL+rPBAQC23HhvARcamY4hSgUimqloommhI6E0g8iLaXThYLl
LbO/Sr6SPsxJraxvNDf2Arrz2SMY0+XntWJN9lybuNt7M+WYVCZjK3m8qMCCaLIO6nvVLE1R5dCl
LQ7ZQpGk3BQjh+vUoPSqMYkuAfpZIKHkSyYM3YyckbdeLroAX/FMgnm6+JCBqU4yMQ1KbelaCX0I
i/hSJNtUJRm+i6vlC8s0ZI07s7IAVaSeh+DLt4DbtTCHPmLbq9bEZhbG3GiyiYLb7Zd8aV4B2u1g
x4cvgN5R7e1D4uNEYilhgj+WrZB+bu97LHSixOLJRJ4fgkQE7CXVQ6qE9ziQRxQ16WSeDyBUy0hX
GYtKrJj1mJOQzHbkF6ttRRi5vhHQj4xwAP/5E0QkzecPPPllwmoeXLkF1PCN8iw7bBwgCetk3nM3
e9wOXEtmuvxb9OXH4ZLPkBq2QhhelYq5goacPEW5s57AlwAtJIvOq4l7xdx8+7dC94a4QVh8qZNh
cEwA6XKOm5pTYYgSU6Agcfonjj7MD5ejLuXHCQ5k4c1ay6wl/ALuMaqdEMa6q03SwyYRO8fc998J
68xBXdcV/ChmanVg0W8dhnW32g3L7wU0mEQZ5buHrHDGs+pZDOBUL49paPsdCoHDoIDSvtFQvwTV
6CvV1YKhRlfwdE8HxjQUCkNvS6+bDR4GD2EEc1Z0uTxL6S5B9tZ+YjPgTVLGmwbE7XeutlBLpWr5
PKay7RpjIway0jIMQJEy7pMi2JeklORTfpoTY56W1VPt+LVbSJZ79TPpIKGggs8+Lmq+KfvADUJJ
mKRcktFTINlH6lm4TW/fOU3J9B3mif4fWuRSGiO4PHrDaZHm6pIfhfME2McJ7B2ymjBP1kL2rs4c
Ho3CNkPIrhcgGsWKVvLkbh77VtmVvnqFqbUZdTqSXx5r5j9rTA3Hmqp682EHlG50ghB/gh2lQQau
pY9w/Njuyuj1AMYCGlhX+buqMEmxnG4WQea5XH/sikMzTvs6f9UrMNBNcFVb8VorbWM0GhgE1Z0O
cHoMIZzNIWmMZMvzIJ0gGKEBdgtl+ER64xzVjugfbqkg+PUzmmcxYjaYDESdWNVJM44WUPfNP24W
3cp6Lb+nQnDrJvBSxI+8x1dUcYvjES612Zwflt0L6MAZYlHW/rUd2H2JESB3zpAg0afGMGmUQbOm
VC+iBF6ZgNEHSnrDPFiASPQ7H7LUjYCmCIo/k8i5SJ3d5baBHrbm3RHZ6rIhodnG4Cc1ETg6kS72
gDFvvfHqlDbOmSO1+klXV0slHUDYA+eo34KbShXQhVijg5LuOhV+gCX4VsaomGmr3deOaUmNXH8U
LmQUEEmB1nRsUDAuFl9QItzY2xERm9TRNmsZ4fm6zVUXpB5oJDk7GgZNo5XMpgiK7RKxMVG94LjJ
GVDygDqFB4RGpYm2Y8YA4sr3fTsyuVfxWQdQrHdjYzlbghWnrgElNebqI3PC0dRgsfzDxIO0CSPq
64HL3t2r3OiSdb379lZssOv33mTTJ8KX9fEa6DiBvIwW7vgXlffNhj9Q2CtyU+GiILyotoGOzCKg
yzp2SCWYuxgQEORy9teQDlyBq4Jjg8AEIOJGI8tqnjfC2HEieKEkNv4BbGzHY2mzLIer/H9G0E61
jzak8UrBdyuqeHWu+moHB5iEsKVaBNffPnzlWIw6bUiEp+lqD0l3G98TgGGz281LMnXgCnKgiwSd
OQPQjaYA2akog+E17yxeGLfeQvHghNFfQBtPGXYqJSNZSMrL+6kzOXW32DZdEvO4ScLOV87SYqhD
R2VsqZelHvIwRA05Y9sNeys/p7dGkwzprrfAGUYeMl+dyjZQcbr94G8LWfldyBKP/hVn0jLRwSXZ
BC7mzwSRBkmPmFF7IKJ6xd8NpcbAQUccIGUnFw31Ji71D5O+0s6yJod2ORsE3cVCoSjWS3Ngwu/z
gQFLkEyCnAa6SQnxPmMCsyoNNVQGdME60F1VRuhVRQk4UTA8XRnjfbriEToiHv1vCGTDgYyp8mDw
A36pKB/gWaYF35h/4b6OrZDEZ1kLw4PrRHdMeIUrgBcGqB2dvhOwJ7ITue3KQzDhtyLcx7hl4rCN
GTMZQLuMVbQTUfSuMASD9czEZxNbgcZuH7WoVmuQCPjSpldTYD792hf6c5v4koT6Xl3foch8NQcl
tBCRV88duAVaKyngs4kAhNiaJ2PohIqecS8I9vyofz0VDj+03kFik3UdggCRabfrm5ojLAlOD6+/
ggxLBcw6KY3bNDEnM3FlfTiIPEbMCIcLIGv+RqAbmKz8pQ0xVgHuTQuolbVhBfJdWsDbUd/LBdgL
LFrGNS+G9XKkd9wERzHq8Puncb7sWiNPyiAN0bcfNApE0pZv9EdNccgoVORm3MPu1kQLt4lHhAt/
sFvZlTcxJsc5TedKRQMShHxe4wUnPmvPwjBO9rIMmeAowsB14uIFMGuojtmA+wS41nrngZbn/ytT
/KA1n8xXzjff8LzWTpoAhF92jpDCNOQYErioVz/kuxHDEIxato82snf/e9TQ5LXRwNDNzQG1Djr4
XSECCIOJHS8DsJh7UIp+w/u7Qv5T2VF8q7qXbnWGIQsti+GeUF4nvGdakV8=
`protect end_protected
