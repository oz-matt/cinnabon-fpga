��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o>0�����Om1��&���5��@egf=�.K�89T�N�4�9��T�w�H���J��{�Ӗ�g�����O��iĉJ����/�}aU���0��.��x��w��}�-��Xd�Ô��m6�|�v�Ush�:��c��f,�4��b:4�u{`'�	�4P��yK�d$��Ě$ip6-�^stz�+�ij����8�?�My���jER4� 
̽mYď�6���*�F~��@�g�n�R��AV٧�q����"�R��:^��4�J��)�����������H�N�{(u�OB�髀iiv8�\�]އ�_��ɶa��y0Hr�ݥ���G[r����g��=�3ٶ�*����q<w%Uf���s��~�k
�3�H���W����
�I��w6U�m��Ǻ����bl�IH�8��
ڱX�'���a<�[[]'	��]p%,$�Z ����Ԍ�q�`��j��u�-��`�+��-���&������x�� �,[lƐ�5����Ŕ$)�&L>�~�R<�p�D���`~C�klO�T��vIMw����n���*l���Ӭ�\�:J�?,��"��C-�eϪg�Ve�R�Q���G�*�@� ��Ĳ[�	�$ #��������l�Y��#�I��kk�W}���۪θ˲(]��LM��s�~�ū�e+��%ri�S��1���)�w�4K9b�N;�-��Mc�{g��I���@`���Z�x��KE��{�ꜜʤ5(�2����+ܓ�Å�卒6��\�^v9�Gҕt��K�b�2��)g�>
4��j�N�p�+����.�n8R�Օ��怟i�:T
�"���_�����?��t>N
.��Õ���m6���ɦ�ڔZ@���!�.dF��@��yS)c[��}u(n9z��Q���R<�o0�i����Rת��^�T��v�{�%��
R`|/�<�ˉd��"�fl�c3<����:��*ҸQne��E��A/	�F��kU����W�]�����:�B��r5�[zcDC���:{�כ}��t�Y�`��M�Zh�@���;*����'�n���A7�v�v�G^v%� �O��q�=�Δ�6@NQ���^��BC����)/#x����"*��h�	0�
O��W�M*iz��+��c:��kn��\�q #α곤����{�@�F.h��rX�8�]�f��|_��Nd������ơ��8�@�7t����e�������2$�����ȃ�ϜH!��,����p�_Y�����fE(�I�C�)ZB֭�cqR�\�J�@�QQh7����&���������EC�N����Ɉ�.�#7ܕ���DV��ö���J��(��28pϿ� V�C��|����jH�p�������	�ߋ���i�+lM�t�'�ƚ�r^[�;cT��}�W�'&�R�8q��-@��$?A�L�d��;� ���$����	 dd��-[4R��a��Wnq��J�t��".��k��<�j�&D��{�m#È�P�[��t#T�6����Yg��%;�i>4�|U���/�)'E"n����5�w�>;�gZ��G�w��\u��N��v��7�������#��q��RmV�P��A��:��* ��{���z�}���ML%�*�	���)$��qL�N�:h&�'y@����c����Qd�Q�n�D��I������^{�T����&�r�![
K-����NVKh�Lz��$mM)����%�׻�X�ϘaBU�L�5n�q(l�\�<�J$M�U0��w�d�ӆ�Uh(��>�i/g�z�R�-0��� <s�K��y��M������oi�z�;���LcW\q?M�k�!�~C��f�[�8�q0�x��Zr�68�A�	�ۆ⏞�]E$�����;Ң�/�"m�k���Im�;Rx-u�#��d�vez��e��n���<bu�鯜GX�ۃ���2��=G�b�
�D�sM��:���~1ȣF�i�xn�gsv�a�ې�n$�($a4�Z$�ڤo��zi�^����/�=�R��G3�?Ӕ$g�Ng��(��E��ޜ�`8��]��1��`� �-�DT�����>ǔj��X������oJ�����K���=��n����Y��Ī,y =v����L�����I,@:�gCA#�o �˩6�c養Y�M�����n8I'���\�ՃF�Bv�:5=�jRϋ6]�o�M�5u��W�`�ҥDX��`�F����)��2�KQ�)W�r��P�:|�Ec�{�Ť�E|�"�5�IM���-���S����;��\�ψOx���Ս?��ưjI�9M�Q���F)E���Z����z�J�BȋQK*� A|XD�`m��7��8�!Q`��Z��fgH��my9�j�t\4���������@�l�2��L^����u]k�VA �� ���w�=s�J�]uP��32�;~�-T!�YؐY]ᄈ�B�e\����**��،7"P_�o��HXO��4��R�MRa��(������D�/����c���b[.ޖ���gN� z����T �W�-����P�
M*�:����鳌��)R�p��#����k&��Vq� ��.y�:{/�j�X�|�c��lM���݊
�WaIj�2�2
�i�i~�]�J�w�>��#3�_s�f:�_~�n=Sӹ�!�	�_1��Fzf�:�J+{|��؞Un%�Lx�j���F9�sOxHt}�E-,{�ae۔r7�����Շ�����[W�X��H<�	�tYP��K�c+���l��G��@~@a)b��'	�F��t'��r����AƝgi^!�x��������O�"BY�r,,$�l�9��K�ql�{f)4�$�k�T�$߆п �6��	
��г����*���W����٩SR��\H��)L����HOI��"�i���Β��W� VL���� gp=39�L,P�|`0���!N����@�cp ߨ������<l����˸8O����������#�>[>�D�"o���KXDD,?E�  8.������(<w��7ᶶil�q��OI��qz��o�Ϋ9 �xf"qޡ`��N�y�Z8\,C��b=��n�����p�����C�n�~C��em],�L�Ox�'�#ɲ+a��Al�C�T�s_�Թ�A��+s9��+�f��y�c�d4"2N�ү�M@�z7Ƌ\ԃ)2�#1���c���DCڔNiA���/3d�xи5��VC��̀ ��]R�g�A��=ZXlzZ�����2ԅ�wA��	����=Mc��{�ў��W#��(N�K��7F]�w�<!Ib���=��K� F3����5�ΉT'<���i Z5�߻���������_{(�c>��m�� +��t潺+��Kf��G(du��PI
|��J���w���﫽-�'@�0�L��7��C�q��2��:�>�W_\,/��%[t_0��ϕ>z�{7T��Q�Ri_j7�4�^:l�,������V}�H�$ۢ<*ͨ;�Ro$cqj�����٦2f4b��5>g펙|X���W�y��K_�����e�D���x$���7�]�|6Q�h�