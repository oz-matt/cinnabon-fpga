-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
KSsdzwBQaElTXW0U1FjMgIViKU871xDgGer3RZMSuXI4KL+UKn4GZGAaSxt/2HKKRlTH/llNM/hl
4RQ3I9nMRLJ4CEAICxtB6aIfi59N/xkH+pEjvadDVrqQysaSn254UXMETXHYV/4zLhXuydd2ZtRd
9vtxILGPSQqx9jswgqgK/wAlV5LFLQU5zznIIk6kArBZIpv62r6Nit7VeFQeMRAxZctlJnprFR7W
BpOZ9IyZ+cV+Y6gilI1pNlP529NqxFg2bYcBqOvR9Gnxt2p0aV63IOrcldJcCCSXA5H6tmLwbO89
uSYnm5/q+U/l8/dCau/qybpKS2pD0s2w1EU8NQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1728)
`protect data_block
A93/l7UgGKy2WE9yDRr+Qp0JWwfMeXIWKlqhmEz80Y2naKW4rXIAzg0AFLtdCjEqRfkw/dDnFqbR
xzpvk8Plhh7gtnYfPCOVRirHC45xYH5MQfwk7ZCZUbfioW0E+pze1otbVAV3P1y+0NJIhmlmgs4b
h/4zInPMR7wiAmVfCXhv7y4WKAd2KjEfLX/pHCo7C9myD2URZSJErBkL9aTTLmIj99rsmijIJCgA
gDCqfahNIYi4DM9DCmAHNyDJ+eKccAgqsb/OyXr316jJ36VktHvOPvvhyQ/nFol9+1nVYM2uUGS4
MOgKuYhzB+bndzcvAVCDy8aW8kSK7JLBrEMI6OjWCHjastJdcxiEQmN/81F5FhMFmDFboxZOk68i
n7NeIlZS2IuvYbU/HJO4CxTAEy37tCmh6OkpNOwv9vT7BYE3dcqhxKI+TWKf54VUXXq3wbv8orRX
nzsRluRSDvQSfFB3Jyu5aAcn4Qnb6z6wdQIQ729LnH01Au7UAQUcZAEN26GQLeWlOeBeanheKBAq
7eUFL9cLvx2CKsyxBRSFjQmjzH6VSMPCyuzZxdpW8sDEPSh7YLF2bQKLXjBCTx17DIFZd9jfNPfz
jglWtH4m3nrf1iLtqtex+omYszEOGB84DlqbilqRD8JPeroK/+ph3Pf3eZURkeFr3e0vQ2b6lDDL
LABsuj+OsLL6q+kkoduLsqBnaSFwUM3woKTOgPQ+5Ryd/ey1UGToQvES5pBeT5nckwoTtX4etrJy
7tIcRhl2LJwFL6BQ28ASzNxJIT0eupyXMoKRhppv22n9GAO9V3YfypT21pAYGtrfaUS/YrVxl06h
g06ezZIOVuMvnVSsYRJ/sljoktA2mH7SHXOGU/lishy/f2YBO1PGmUmjCNJK67coyH3ObuFeY+4M
EeODHtaKOlO9MhCwYS9weJgY2Cs1fluJ0d1beciqKOSUlumaC+MiQM/JVT1k0zGO7Nxy/vF+gF3T
OJknRJ3I9V/AOlFAt1EhWO2lV5zoB5XbXKJ0REcCUVgCn18qXnDK31icu2JhPK+cDfgIfyC461rs
b0vnEDQ+BmhXd4Cry2HIuZwP3X83FH8lWHUyWnjEvb1xPWxGnyvcjr45yzSXRvANG2ZHJrKMc1h/
TR+m+AVgA8na9yorRI+lO/G0DZ/wIW+RhFEn2KacLk2kLJxabj8+cQtAoINJ3EU2MegJu/07i0ii
ctwpJ0zx0JoisVLi+7V2phsySwnRVnRIzeJfP+Ve0WvYORE5n4Wq4v0X0mb3yzE+C5ySm93rXX2q
/iY/UqO8bfHOsyivSgRnEH2CNJZVe6IuMp0fAE1uqcwmP/6iGpROl1ku8etcCR9vDOFFjGZJStiV
8gWVZrkReLQmK9EZimt3NXHAM0Mf0JlaW2ODbB181BoRjQhZS/61eDRMHMQOaaRns9b56SWUez6v
S4iHzeL3qWyzqjp3OV9Yn0LS67qwYbADSImY4ngSTcFH1xKpcckrWjCbpmhQH+U3lE1vCS444Bei
YBk0Am9IYMoNflXpwahoKmaSfLaABumFDtqxX3a+gOb6bH6Ei5PvIfbpwKK7s4MJobiUDa5A/lal
y8iYhXvnByBbWQssxcpNF4X5M7jlrTBlUBAxz3i/bnlx8AgPSTorkodUAThpOjAS+Svy3geFFS1c
84TFohv2t1Yk6x/7Qv5AEawRukUFdBB4U9ViNSXojvlD5M+6KUZfMXFSUl7G1ryPIyRT55OcBXVP
5OjBgEfnBIzZcBvfpEJSmTCxehLL0v+LXApTjnTpczvCeOtbz2HjQdZ17UPETdVD2k447OjZkWYT
T8ya3uH0H+HFEGfneBs0g0goymaZqIVJq69Fqt752u6sUuwQsafo2C51JpuTW04YZdNNwGiArY2Z
VgFPCWYpjXEioZOTx/dEZAlZBSJjsxZxlZp78Al7jxKs6RelJAtsO71c6E2JxILhWgeC6OIRCVb+
D0JiHHfu/NbEyYA6Dejo98lEN85bIefFVIWovO76oGTOWxLtd9LP1nkjSrR9fVj0SX6CpzLmKssQ
teE6xje8BjcuSeNCha/vZ7YDxNmrwtonibS/pYBszJbiz0Rz8BPwnWbLISWXRakyCIH/cqbgcxrA
590oJmG5EPTQux3lXQv15QIaiZsHUxgVjXrsULrKeFtbZfvIrEka7DTrWaZkPrK9vw1Y4SNOe3ib
nG+P9QJknu0nSthPZIqag3z5oYJ3x49bc/qyV+27drd7QTgwWTxVZF7NnfW/OiPNNeAPgEsX0o8N
xR9TmWw0AJrffaj4M6g98G61
`protect end_protected
