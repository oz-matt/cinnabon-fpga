��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o�'�k�l�A�.]
���He|���(��n�0�:v�Ziڍj��E.�Gk�i���QolR~�'ըD /�x���f&o�Η���`M,���f��8Mb�$���F-i�IVz�i�~Lh�� ��r?���.ot��ea������,�/@B��7Rk)^�x�T�]�MYh�Pba��Ug.���li�唉���#-��XR�Y�ڇ�������Ya����:��8�#y��+���=+��F>�Qʯ&���7���鈗H�޼/8�t����5D��y���$M<�t��U�/�?:�+�>��n�QPe�_��;�}0+�ZR���\���W�P���BLHg���|g��]
�#��}ޝX����E�F0ѓ��]�_]D��=�C9t�P0�;�X�`��Du�I3����)�\p���]tnq�[�d�X���'X��~��Yzw`-�f�q��5�W-��dTf����o�[\A<����]�0��m����hx�X>tZ�$?��I�8�A�t0Į���X�7�����P�������q�[�t�Lv��4U�nOR�3nCQ
K�M5U��WZh,J�B�F8��6�i����,�*��|X9��
���m��*r���ʧz�j�̃��=q��@��
^�I�~�H-��ш$�+Q�x±���n �x�Ջ;�@ �珆�����X�w�_�A���{u�d/\��5��� ��t��&xԔO)�R =L����2��K�� �X�O�S\�ƪ�E�rڧ��1
N�D�0��a�պe�.3f]�7��� ��cF���b��+0�B�Z:q彎Y�`u#���p�OT�
���qF5��/�]�ʢ �A�,��Q��rc	�I��.���$|E����w�.�PX9�#�L�X� �N��I�E��Ur�������]F�f�%����^*<�aF��b����b5lk�E�� K����[W���چ��R!�I'�_#O_�_�#��I.TY�Ԧ�������U��Ɔ��l����`����NJ<>*�YE��)�%[�G�\��n��&�pk��ϲ��k��VN�8���(Csxl۠'��Z�W�	�S��'[LR��GhX��P=>JN;������a��ΪT�dY����-�� �S�ѯ���ʞ��T�4�Fd	�X��<?c��u[�{��K�3��������&�pd������H���K�j�籩�mi����M���3Mv�皱�{�s?co	?��_���IAf���b�x���,�gW1����0�eL����K!f�h��p:1N�G ȣ~�5��Y�˚A�\o�G �9�V5��|�^u��p_G@��<S�fd}�l�#�;��j�ZQTS5i2D{�[f���Y>�Z��۩���_�ݔ,G�W1�9c�� Bx���'b>ڞ?��à�T��1b���l�)g���#��AU��8�ѾgS��{A�=�;R4KX��P˳f6�ĩI����vE-����u���e��$<��x�+��iQcɖ���/f�g{,D��^��	O�x\?K$l,����t������P^g���[m�q�[&	�����2B�����o^}�iC�5x�x���;�����g��}�T�X�?�,g�D�b��EǾ-�X6�OH` -�l��ڈ֤��/>wPzg�|^�r�9y�I6��ۺ�:vī�]^>6)�84M��B�Rck�zIô'-mЕ�n��C��P�Ut�}��%:'c$e����2�3<(m�m��vhwr4uJ�a�������,�>;\oX��oC�!�a�N��U�à��\b�����@�����k�
��o"�p6�)y��zPR���I�&�4�'��R'�_��-�̑;���P�?cwȅ6?��ga��*�pD�Ǘ��i�L���Bt�Ȍ��N26yN����滆�ڻ���w����n{dS�������K������lA����ؕ��6M�t�Q�[9EK�E���C��&K�Ѯ��TMO4]/,+K
��=T���yC��!�:�Is��ińu�Q�6"#؈|����}��s��a�1T��
�
���$��ޝ�T��R��5<��{)�H����K䤁bp io�T9ߊ�&�ǞA�}�R�F�R�m�CN�'˄7�Yk�Tޒ������Z\;�Ts�Յ@a�9�Z�.fc1�����T=�1�8� �4�S_?�CþIh?�khs�1u�l��c����[
�"?�.���@�g��fȷ�m9|�v�������h���F�lt��z$~��!bC:z��״.a@;A�3�}�o�gwZ7M��F7#�[I����\��Z�18l��ta�1�c~���y�f�b �E�Z�O;\��P�*��}M�>���� �������S�����*��{zo�q�
��Ni���#�[�����خa�J�����ĳ?|��A�op�T�z{���jb.(���S��"��^�~U2[�Ð)񜞓f���sɎ*�e#�EFQlRBO	mT➩���a��^�
���`:z�,��}ӳ�s�R}�K#�U(�	=S\����}*�`����i|ڞs��q�+%�U����G~��	,q�ۊ�BΟ|�
6[�0�o�(���ҍ��L�\������D]w�h>���o���أRr�Q�25�b�᭕\�)��Y!�S��)�i_�?����W��^��3JrM�*(>�gf�uH<܈�iJJ�T�)�H�����[�m��{%�Q���a�g��|��G/���Y�a3��px��:R�e��Rb�#QᾛF|�V�O
8���Rϔ�M�ό[�>>�ZH6r�j�WJl����mi��� �?��� *�e^�LFb�d��H�n=�v���ҥ�M`a0�c�T�3}����;n�	:�����E���Z������o�ڒp;Ԡ0��e��s��\���Ʌ%%������aV�T��AYP��� q�y&���(�W&H�c�[�ZT��c�R�Bb���3v�������"��Ē��U��'^�$ȍ�!�XU�,��|c[������!>��=��7o�S׬R0�C�Y�1(%���T���fQ34�G��ص^��/���0D
h)�z��.����H=����w���a�U^؋��'���GvT�3Td\ss�/�}.��?�p�:�������-�����aI�h%gI�ƫ��0�9�i.�o�O��y��_��rtU� L�w
czw�=�Qv"���jd�Z
��������.1Y�99����eR�ܚ��W��؉� SO�gɋ�ZWe%�����y�:�W �U����I�U�-��FP�C=�ѭ��-J��N`���Bv6]	��"���y��9�iN�VD��e>Tk��C��d�"���I�G[�m�D�dg�TZ��@/��a� �/͑0��/��Fh�ǆML=��Kv���k���?�ժ���_�ϳГ\����$v����i�B�9���� 	��k�4����3��_ډǙ<Z��qie�Q��p̫���+���<�5Ru�ϴ�W����"%4y��ݷ���F��V�NE	'F��s��Ql�~.v_�Ň��Y���L~�xМ�[��B���{7q���%����xf�:&K�G��L�ِ��ޕ�3�Ź�6v��N��W��-wf��3V���s��rW�O:��q��L�:��"�ym��2'�K� ^F� ��t��'L�!�e��2����h"�9ʠPP��۸u��P�`�:id�8S�����\Hk��~@�)���>·�p���ӻ���|��aTp_L�> �O����肾x�1}r6�v?��4��-��aQ� �����<�U�L.��+,��n�y��G�0�#�P�6�c]����wuN|�����x���qw��1��7r,��^fdz{�=��èT�G��)6vA�`%ƈ��ɪ�뭶F��b:!����
b�������E�_� @:ڌ�!��t���N�>˗��A��B�JTc�o�z,����X��t?���, �b_��vt��Y�S;I�#$�~u	� ����*cb��6O>@~�TZ��<����\�d&��ly�5��%�Rma��v��l��Y�}��J"j�#|֯(��F՟��QqA�ǥ��b�d
�VjAnˆ�El�Zm&��5�T�7�ȧ<�U�=I�4��iD�������������T�)�k�'}gO�p���Mq�Ϯ:�{c?oKM:�3T�d��N��4n�N۫�٤X;���#��J�� C�GvJ- :�T&�R2��@1<�C��ew 6��U���5,�͆4�.#���#��(�P�z�$i�T���H�n��E(Ύ�p��j�;oh�U�i�ŀ]ӿ��/�q	�}A��7�{+m��OVڹq���C-A8p�1�b�o���/-��<��|A��Ʈ�wZ&E��kGr_�X���'�O	�P<��06�>�r�l�N\�=��ϳ��c�8��*�ݳ	��E�?��������M���Udq3����Cn��6:�N�>+b��&M��9��050�Q+o���x��G��׃���ZE /�u�bV�r�����y>B��fb�R0��wcc\����?����L8�!��r��ѥ��.�
�z��CB^�!A�	m�x�fy�?���d/ ��o۷ ������ӿ�-�"=�e�f�7l�A������_��/��T������:�[ˤYx]�����qE~� �Nn�
�����ϧ�х.˫;��P�4�/e�?F�u��P�S��
��ʃ��|����	?�U�����q��Nf��8(�u��S`��TyRƍ,�h�s��E�b$	ځ�g4ݗq&1��+��@�LC�f5kw�ʫ)��P��� �&��Y}9?;���N�WV��M��Hz��5gݱ��b����c�D�*UI�9��v0}H���7ٲ�Vys٫"��s}�P!�����)���sȣKZ���|J�R-��J��� ��T"�!�B��ʮ]���Yڲ�1z�Ax�X{����<_ؾ}�4��t7=N��FI`����5�z��W�?�zp��$�gao�60����K�_#�+�T����m�K:���ٷ3ܔͪs)#����ui�9�� h��1 ��*F��h�^r��l�[��U�B��#�E�4�dbݞ�+�V��&��Y�}�]׎���tl�T��Wk�ʃ1?��/���瘃�MW@�>�͟�*��*/ƍ�ەl�d�}0\��&��1��'{G��d��#�s_�kMa����c���4�z+U��C��<�ެ["O��%��4�"��^�,��qX� ��a`��<ӓ���:�w�N1s��	�Ș���A�4eƊ��7y6u�Ȕ�

��BiD���k|�RO�|=�h�So�oP5��Ͻq�<�>h�DE��ܥS����e�e�?�dS%5�7p�6�,�\R,��r�Q�>g����aw��8"��p���I!.��T�	�6�����ꁏB���"�f�U�Cr��"��{�k=Y��g�FS�+�""�/��ZK��û�n��[�3y�;7�h�l/&[tc�$�CO���a���,�t�s��l��(~9F���7vs�#WC �a�Χ���٠��#l/蟸Bi~Ҩ ���1����N�t/(���5���,*��ś��+�^s��q�����Vb�s�w��Yk[P(������?i�������t��f��S�$���%��+((�b���#凄r��[!��P��mM��x{��_rW�č�4��S����̘T�a�a�#Nl�:�6��{g7U�����6��G;��&��Љ�N�Vדm�ù�X��tYR�"�OW[n�QB�����i>����1($}B�WNO�o\Z���N������Ĝ��xc@"�p�$\�ΕoA�6�\��e[�#	�0X@Fs9X��]�����z�V�3���<�Wt:SB/��d+�Lr��긂�`;��fs�qT�Dr�n3Y�ԅ��";�c��q�^y0G����������~��cgTLQV�IE+/��.��|<\F��(�N=����|��^Wf?Y���N�Y{��"¤��GkXVT%��4H$��%E�� �����JE�E�O��롗���1�|�v$��VS���O�~��)YÎ5Q�OX�E����� �Ȗ�L(��+I��R��x�	7�DPE!�-���T[�%� ��5�e���i�v�Ed�`�";������.����#��yƙ�'��@��̬���2B#���귈�,
1'�A�&Ԡ�%~Ɍҩ�rd*f�k�.�L����p\j!�S8�AY^B	C��^��ڟ>������C8�`i����-k+��lwx?{��'��a�xs���L��cK,�-c��y�A(t�1�{LcM��0̽�������H�Q"�F�9����R�2�r �� ��ٹ,|5U�ηP�.2gH3�3t��e:'٢mS:2!֌�'��v�-NN��[0��{����MOt�G��4���v�p���$�8O5�(�Hc�a�g�E�WS���8����ѽ8-���0Q�p&ίc��P��8b2C'Q�螚~��-an��%A�g>Vk��9�D��.Y#�R"�����}bp����$g�tY��J=5��n,�Jtzȃ�N�:y5
�ǖ99L�,������%6��}~�А05�5�ت;/����[��?��\���}�xSϸ|��+:�>1�9��nq+-�z�58/!޶��-�F$� �ܼ�<� �{�/�g�2m��7k:��i���׳�X��/^���ɟ	U�1�FA�TLؚ�wW�5%Y� [\\��B0Ye0jӆ���'�1?�7�� 9�C��2�+��xQ�)��6s�e!j "'�0�2���\������3!�)��f�]�n�#�=� �i)r5�3�s>O��
���!��Z��G���ݯ\�Ფ������?�¯�T�����|	70��C�Wg�[�&��Ŏ�u����q�T�H� �#9#<X%�.V�j���Ka��l�տ�o�ζzR�#
�<b4�Bc��5��?�b�v���ֲgA+N���+�@,7�,cl���y���C�:�|���k�K��/���*.����z��Q�W{i���4���C�/��Ԝ�{�+�.K{�=��J��U�3�N6�Ⱥu�	�3~�ƥ�J��V���BքA�~�����%���AD�1��  �L��*x&�uş��Gl���s�٦P��Y;Dj�o�d��������X�  ��H�0�9�V��w� ˩���)1����7��	�1{���J��b��㌢�ДU��K���T��B]�s�5N]�uX���p@u���K�4^3횔I��Zʲ�(��(�}5��\I���K� g���&�/D��L:9�� �)t�Fzu�'k��ma@��n���)H�Ɇ%�CQ<��7�j�d�?&�R�p
8΀�Wz0q��{M��۰B��s�-m��y �b�p�R����%2��&��*mO_��8^�`߱L��ꍬ�Ĕ\?<���،��1ַ�ߢ'ywBG8���4��i]���Y�G&���ty�J�W�@0Ÿ*H��{�5��V�����c���4r;]҉�Q��w8O��Y�Z�&��"��D%n�~=�����\�8�x�e+�Tu�P����_�0����4ߞ�jȧ.�G�T`n2��V0�\6�v �m�?��Y¯�v�2�Ͼ��A"������ǻR��^�����p0*"|+z钒�8�P��!QkA����f	�S�j�
[��j�iYL���r�ܰ����SJ����+�����Ѧ�r�W�ƩP��	
�7���Έ�ɂއ~㲬��w�}�V7�����
�������q_4������a��EAXP�ϽR�x�p�R��FfH*���t�rS��c��z�?����x���KѨf��D��}�	�[JK6��o���o�kR)��Ү�ȪI��b"����{
{��;��s��gL��Q��R����^? �-��g)?���_�Hl'@����Q�m��o�'	k��P^Se�U�J��L3�mg� R^��u�z�l��Fa�G�7�V�m�[~��������и��*�U˼�ā�>�_�&�7U�@�֬�����]�Q-9��s�^�S�ݩ?�Q����@��}����n�/FI�2��r8��������L�C��Je=�b��K�j&��p�D�Ӏ��F`��nm듷q>N�\����-B;��=y�b҄��B��G�)r�T.��������x����Vfq��!D����>��y=Y����;�1s|��	�����\�NBhUt�<]�c���qN���c@�C��cZ�K�sq�����;gy�f�O��!мC��\�y���XVa���F�|�g��ܾQ��Un�Oj�-��\IX�8��	(#�)�o{s�5�>�Ʊ�SM^땤�
z����$߅�9D	�p���ڃ�t��1�@ \�F�ϰj���8���!-��^�Ҭ��]C�g��?
:�U���b�vf�b�,I?����Ƴr 2�ㆥW.[3���R2����:�(y�+�O�!��x����/��S��J�O���ǉ�|�����\�%L�
�[~��}���˵�J%+��p���H��	\��p����	i��fNfa�Z�o�$���iF�4?l�1OM����BK59+,b��O�/��_����s}r�o���7���?�>�C/uȇ�L�%��W��w�&�'�kh�e&j��G�q���M��2wu�6�x����d`L����f��W�z�7�Qa'���/���AH���4�gPq5pb��a��Q[��A�^���\J�.ޯ�)�p�v�u��`�������%���3�O�Tݴs�l���>�:1L!�8m����񞬁8JGU�s���k��?k/��5�{�V���5�A�S?���s��'�P�H��I�n��G6t��mlCq&��-����׈z�h'�}0�c%�K_h�۵�Vص+i`Capx���\��|���H�fZ���܍�r�����)<�� ͠#�S�n�\���R����R/�oY/c	tdZ >	��9��=�:�w_���l);zQ�a����!X+\C<L-�GPD�lZsO��{WM#f�I�?;��� �xʈH�pl�mS���٭?�^���\Զ��� �<͌���*3��b�S�1������kXb]��xG���̱�c�	���#!���Gȓx����{�:͆O�杓��n=n�Է*L@NDQ0e�a���m�̧H�Y�+��'��p-EcEр��,���9m�j�Yt��-� *�+�r�:�,�_��=}�,��9w)�m���U@6�'��\,�	[�p�8$�|��59�Y�Y��9c.F�e7Ui����UӮ���ـ8��>D:f�H�����A��zp2���D�$����_@�Fl	�3l!����__Q���B#���{}Ȃ�#�";U��z�7c��Y���R����V�F��ǆcS�)h����ni'�3�<��Ŝ�#H���xd,H%���C?E%eco��K\���K�Ȩ��h�a3	�@ �B^a��O�뀩�(y{�@�Ԧ.����C�v�=�n_��f�V���3�1r~uw���D9S���"���o�N�p��׮:�	S8����-��T������
��9S<iG���wy,s���0������z1��~2��d7H��e�RX�·�-G3A��4+�
I���{BX�R��m~��M�!�9B�� =M��}��f�^�ރ#E��g�aܖ+PK�� �x������^�q8���#mr��o���q���jg��<�l���<�f+�[�zm9�"\2(�	��Q���ٌb���F�Ŏf��j��_]���q�<�o}���2�9BH�e^��Vg��9����b��^� |�&�x=����4��4�4N��{G�%+�2���E��
�E���i���/��ĺi��79*��n��x#��Xr6�=hoHL<$	@K�Y�]h�>.�P!>GsƪM��Y��};���X:
_�5�;y^']�݄�Z ��1Z�{��qxF��pv�4fm6�,��#{�3���+S�p*��%bt��/�;u�{�xj�Y�e1�x���f�Ċ1B׼�"��~��Qx�R�� ����*���VJ���:{�r�z�5��� C���օ�Z�ߴ�;9��y��^˟�r��u"��a�jsݹ }���ꖓ��'����y��&�)nm���"8�� �5/�� ����|r�Y9��
C.R���X��Y�g��������ꭰ����e�����oW"ىY�clgB�/c!a��E6�q\E�V.����AwA��?Uh7;��CJ�0�?����w������#������^�����{�{�C��ZN#'{H��0��}�1�>������Lk�[�,����!]H<���r�S#�[a�2$m��\�3U�������8������A$ϥ��box���U�#\#8�X۟0���%.��m�lX�<��;{ǏV�����/��3�����\^.!�ޮ�0}CNdM�2�p�i�p{�'5ħ;��r?}w}������0/K�BJ'����s8�sj;���h�*��j)b]�X|e7]�I��:J���R]�M*?����G�S�{G��[�m$=�t�y�i��
��ʦ�J'��d��^In'����Lfl��85dP�A��{�}i���\q�~pE�)�z�f-���!�#j���r�̸}���{���@З=� ��������K��?��7k�TXW���M�A�a?�%僌OI���O,���m��q�����"f�?�s��TLb�:Y:�^$�*,6��ã����m�2�-�j����@�`�.L 1T������(�w�]M����Hsm'���ٕ�98X����+�����M���̲��U���&�49��3,o�^(�[��aBo���,e��U�f�$$̸� ��4���A-�e�;�Ɓb(�d��O����q�����f���D���⫫�>V�:���"��'K�Uf2(I��9#װn����}qL�����̓r�f\���i�_�	t������ya83g����V~���K��;����^l|���w�?�C��&��DиW2��.�H��xmo%^�	�z��T\�HT�Wl�A�d}ŭ=�Rt���8�ծ���	h�i�cF�R�1��3zזO��ܺ�I���R���b��I�9s��,���aDP�'ZG����ς&a�V�� n��������>�I0�I����ֹU��"P�x3R�	�OK��!����#nS��`B�k�j��Y��.���S����Fy�)�I$�(K�}@��g �O|a�r�A���?�����9̈��I���µ�ܙ̧�� $8�>��,��ma�K'W�x�����W�i��1�u_�\Kp�%�o�4�ٍ�&fgώ�;�f���Si �xiZ��%��T/nf�����̰j�tL�%sF�������1�'u@ �MP
h�5�/����{=����Tƃ7��A��_h{/�}�+�OU^OR]lWݛ�OSNb5ED��'>#/Mm��L��SPD�A{?c����8�d��Ѿ0E���Uj�UMPXL���=r�&�s/*�wf���%u#����;
qIo�?T�aO�I4��财��y��j+@��\�f��:�0
#����I�g����g����iۦ�%��]KGׯ���3o��F��g8O+���~���~{@�it
��7�p���X҈�ds&ꁣ�H��hZu��n�D���o����V��Yf�c�A�r�t�1/&�����)l4?�KYx��K�+�MA8|װ��U����Cz.��L��?��8���r�5٬Y��Y�-��VY�z�ϧ��~Ot`����9u#�~�$����3p�X�_q�H�U-�8	:)	bc\j!�a�"sBA
]�`>�Ia�X����*uW������F���̾H�+P��Jݩ�\�+˂^v�Ǻ�"k�J6�/��W�7�;䛵�kP�!��PHp�n�*�����$h���/SA�RP��� �o��>д���j�[P�6��s��͎E����Y"l>�w�?���L`�#��F큃 �oܘ�<�n�@����1j�;���Pm_q��
_�� ���N5��6�%LF�����-��!���ORG��F�~_D�Y+o]�7[&�CI���AB�,$�a�����W�Ԭ�����(=3��v�&�s\���-I�IvC�a��ΆL�7JK\�	���������lJ)}����ބUغ�S���BUS�a�Pe�e�[������/ �"0�/��j���AӲ,�W���S��������vGr]���i��)�e*��4i:^�A<:.���sQ|T�'"�d�$��2Ƶ=�zN�	lA�L{!���2ys+�a/��2������6�������q�����k	ߨ_l�&ܒ�Ӂ0�3����斠633��L_�����D3�x\����H6�^���k |��>�N�� ���*��Ùn��[:bVר����2�\�θht)���,����eۙ�\�0�;0���Q��k4V��b;�҇[���D ��h5[���(c��X���7������'G�5���3���@x �ԍ$�����:�� �E�o�>�5����
�v�l螙..w�>/��5����	�6�I�f�HP#Ε��}�����&��x���v�V� �g��IN&�G���Te,�d)?���)���/r�F�s�*&f�Δ0oc%4�N��Ȗ��
�IF�cq\������ɄR���T�F�ae` ���s�|����sU�����w��a_��K��M�#�h�@�F5�R�4�ul��<��5�z�!�=��íWbi�ͫ���x�JD���<'��'���-��F�:�[qY�K�@�]���X��J��޿o��w�y�nG��(��'&��vr�J�ZY���IⰣ2���]�G�����.�$4pᓶ|dɝ֦�K󊍃0V�
m�T��yڀJ .�v�ފI�����:`����0"[F�'�Fg:�%6kq����G�v<�L�K�!��"���瑄�h�¤�S�m�Q:�ZH|�s�	���rQ��r#؏�zC����a!׽l}�ӕ~�t�T�[�v�hǾ����T㮟WB��F���MԬw:q�U����!B|=~�15�5�$�m=�̯����JAW�|"CAhOyx�������*����H��57Ra�\n�����(������Z���ɱ�>����@��a�r�C	%.��M�@��L��2��w*���)�Q������v�j!2y��q6ш"Im'AK)���\G�{��AV��?#����S�p�]�ۚm
�i����E{2Siq��ZJ̔v��^���>���E�Bg]F��*dO|�X�1��;e7R�r?��ot�Y�Y;�k�y���v����(�D�(s>��ڢvX[��`�� �|�ɇJ4�չ�v�ɜ3�L1����6�0w�@kGNS��]��Nt�3y8ؠ�Mo~U�:M�m�/�'��?n�V��20�y'��>m��nԤY�fr�������+o٩�h�o�{��)�Nv�cQ2�¥�#B�37D�塩��u@ϷY�����8f�x��T�4%>W޷r��^b���F�HU�y<o=���`n`�xԸB�͉D>����C�oYy��k�Y���E��ky'08�	���I4/w�HǬ#}UYt2�"O��Y�hS�tƍ����3.IaAo�(C��V�<H
/#f?����3 �u�(�U@��!<��"��N�Jr��>�S4~��D��w�JÏ�:I�������	X&�R����Ţ��b��y'۩�Q��
ؽɲ�ᱯ el�RDܿ��H4g⡾ai�2ɹ�!O�w�*w[��1�<�By�*�s�����8�i]�%���8�~�~~�)2$���ӳ��6C�~�g��-��)��J�l�Z}_�8���A+��^�12�rǜ�hJI���#	UՏ�#~��)�T��\5zGh3����u�]�ܢ��\9CUyb^<*�i�a�p'k~���s����3���A4j2����&���8a�#��=�IU{g������J@��q�q+�q�Pz����-6���j7(�7�6�}�ѳ�����x|��h��󣬲�UDL�Tk��I��9��r�WTIJ��͸v&+��_&���z�z�\3Ɋ2���Z�Ŝ9C�[:���
�>#����^l��G��� ��H���V���S^�ژ�V���;C��� �2�գ��z4�3���3i�����ڲ� h��J��ʄ�=���f��k��y�����)@�a�r{�k�v���	[wn+f�/zI6p�r2а����
�2�o9�{�J��E����FB���3�5�<���G_?Q�y%l��� kCw�Ю���z,�����{���p�.(����<����f8��W�W��q�����0�	ұ}s�� %Z�OTD.�V��_�R��]h������90y�xoމ��D��	6k8���$@�5�F���T=�e�z����mY	��6�ޥ#�a6�L0����!�{6�u�DM��Q�n��~�tS�TR�$}� �ɣ�Z�Fs���ݟK���DO�!<Ԅ�t\��w<N��� �S�i����\&]�-,��M��<��z�ocCY$%=
�u�X��ҽ��.�f�br��t�ڤ�gf�ݢ��9��T=Q�<�0�|K��
��m���/NᾣX��)��뤏�Ih�'>)��s�.6��;������Q�Ɗ#��WäH�'�B��5b����`��g4��<��b�~槼�I>���kt��^`��(�-D�#� &*�8�Ef���Ȉ�N��n5��B�D
H��7������S�96([:'���fk��	(H7$���OAt�{��AE�����w��P�����X���{�>Ɩ�����nI�)����$�!���k8&P�;�u�����[�q�L����n�qAnJ3�H��ۚ�����G��Yh���ܵ�(<N"~g�*�?� j���uSԌ{[�`K���p.b4����)�Ŝ������]P^}�z�`b5�yF���}�U��/+Q\��6Օfo����̬n�H��ML�g	����X'�]�.��5V�"^�U�\C�w�۩�I�����h֋ 
��mõhi]��d�$�)gUI�Ó!o���Tyn�0N�}3|f����/�#t��|{�<`��$d`�I���m!k?(7ĸɍ'��k~U7d A3�E�tݞp ��j^���QI;y Hp٫Pg�e���٬=_�ڨ��6$z��x��R��'X��6���fڒ`��*�ս��#A��H�8eBZm�o���t�/=N��g��`�P3�*L�q�$S�vc���{�O�Č��0e>L������:���&Bj�.tR�LF�slqlVh�Y����`؏ͨ^h�3^���ڈ^غ��Ca���s����?��n�6;�.FUg�>|7�mI�y�g� ��ZG�T��I���W��[0g,r��A)�ލ�S]QI'��(R�֣I�!�a�
Ga�޴C�IH��j�wآx'�m���7���V�?e-Ӣ<�j���:�'kv!��B�Ip~9Q�T嫘�* @�;�����k^�Ψ�P+���󳴪6��'�D��`�����6�,�+N{E2��gפ��A��R�J�Z.���*
�<��]���dpO4�C�k�����+�5+�5��3�qw7�-�w�����4��B�DP���������{�D���a�OE��JW�>�;���G �{o���G��a�%P�C�lf[Ha�/�̵ʰ"����q�qzxOf,��|�eZ���X$rbFݣ7v<��Ī����N������1��4�ZU�:�!�)/�B�{��{s}��#b��>�䰻�)�=�)��ȋ�LJ(��1�v�|o�J6�-�%���塚�h��2�<���3l:lUJ] 0B�:��Ȣ>5�1�5�Wwў��9Ɋ`�h=,
gT�',J�iV�60�2�e�K#���
2lj����N�T��yR��-�/}s1@�p�%%�<����C2�0�'c�Uݒ	>CD�9'�b�M�0BkB�?V�F���91��R���o�����q��lꋝ|�m�x-�g��KogY*�J�OU�ʚl��$ F��z�iC���a�[�p��H�	9��!gI����}HϞa�W�f�+~�Su	����j%op:���s��Ƕ�X�%W�"�̄�>�/��(��,������b�C���2p/��?[��	._���c;8g�>{GL9W3�l�����T���L�l鉿�O֕����ڻg��}n�@�9��18Z(�H�:�%;b	�!B��������`���t��+�J�6,��R��7韚��!��
+�1��Č=}v-<gER��M�������$��Pl|����0�B>�ɸ�/��y��TD#������e����r�Kɣi���+a��k�ԛ����e[���a�Z��_��0|[�ˀh�����"JlA)WJ��'�|f"�g���0�$�Kb}jq(�T��̛�
9�ӻ��9-�� �Pr����O�1:r��Ů��:8*� 3���j֖��}��\��&ץ���yO4;� ��{�M^杏����+'�2��-��Q���Q��/!��N�t��b8C�'�a]�����.� &��F{��Z��@��~�#��M���� �^�	O$cj��}L�����d-5����7��w��H�f���HC�`ꋧ�]�X��҅1�ͨ�Z�C