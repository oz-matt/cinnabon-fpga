��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&oi쵋OZC����z��"���jt��M!\�T��x��gg�)�s��&_z�y�=N���|<dW�]�E��'���_�p0���'���eN�]W/���bD�r-�*���,��6�*G?\/�SF6�`�O��ys�h?n�I����>q���3��r5�����va�µw32�;�m��L�
����@G�骥�+y�6�i��f�^�uK��!��G��[kP�.�V��s��1^�Q�仕�,+Jv�K����x��!啳;���S:8�ؤ��6��q�R�NaW9 v�)ԕ��sa
~���癭��1x��#_���<�ۛ2ʽp����)�;��G�P����N �@LO܈t컬.�9x�A�z[��+Б�(�}��ۏ8��X_r|�̍���3����iFh���b�,p0802�����U�X�?_֗�Տ�z���;��V6v�ĩ�pC�2D����n �H񅺿�P�a�j�ᷰn_�`�pe��4��	��%��ݜ��Ԋ�5�ܠ���:]���?F���S�Fu	��K��\j�O��ԗ��:ֱ;���Y�������ﵜLb�/����S�X�ɴ�VoP_���{�v�e1����B�Z8�*Cd�GY'��ђ��`[X�5�s��`�q��{�~���Z�}˶�q�>-nV� �[ʨ��SA����GE"��'L����p+xB��Շ��k��Fe��ʏt/�q�'F��k�C�dK%Մ}G�o�>�P��(t�{�����*=�6q�X�s$�AzQ�q��Dl2y5���|5�j�T'J����uY��k[�+��&����ߑv=�w/d�^4LR�a�aiL(�6=l�>�9o��zX��ݐ�]����^�}P���	�M��K.�.m��d�א�x?̟�em��܎G,c;��l;nY�kC���`��N�xB4/�nVsL*���O�Z@jR��t��cT��d�
WJ­B�Gc��)G� ��K���Y���<)�95��� �38`)�k3���y�[,�^Lؙ��5v��VrM��_Yyq�?̍�n٬d�N�A����zZ"�B/�O��ڌ\�h��a?l���xPy�Wc/��C|Sh�Th��Pw�Q��C@����](�<Ue2Z�G����c�r?�q�W�IW�Q�����";n�p��ЏW3���L���$R"�E��$�����6Bt�\��j�����A!}'P,aB��� ��\�zP���iē�?8U�$��'�c�K{y�OiS���W)���vG��ʖ(�ڐ; ��k��*6K����r1�A-�_����rq���%���_�6be@>s=��<�d���eXJ��݉Wi�,�i�j:���/�g�ok�}�}��!>�WGAbį���Dו2�8���e�N��6��"�s�E��}'��rN��c^������2��9����Ao��9��"���������Kng�>���>i���UˑF��I�+��@-���Sq�vŰ�/��J��{�?��̟�����Mb��C�B�W�U�R]6 �0	JWqyo=����Qu�]���1��-O~=�^B�����:D�3�S-(N����`BhG����s�P~�V%}G)d�7M`�C	�XƲ�"�ƥ�&{�-۸c5:�`"i�fSxy)[+�l�J�[a؃J䌾8�n��3zשBC�ԝ����.���Q���|���-������)M�V<=�,~���룕b�1�T)�Gq�Ɉm��c[���Z��Ao�<�Fœy�ssꭐ��?T��W٨:^�>��|��B�Z
���'�Z��Ja���D�P�<th\��`���ʵX���b�u����֞��CJ�P��΀���"�����#�v!8�����5{��>�Iݕp*vQfD#g�`a���/��ًƘ���������@x&�� ���	u�{���P�h�p�im������C�Q�2嚭�Dk�nVݧ�h�$�����G���s_�;��+F�-մ�a�D �:؋�t���܋�$@�U��t�T�I�e>��$(
x6kίX�z�2��^��B<`Χ�[�e ̓YD�BB�5����m%\�'�A0�̜���Z��a<� i"���@�n����%wr�o;,Ey���lhr�g��x�m-ˢ%I�{��.�7��r)<��|i8

(��P�$��p(���׻�ͯhv9<j��kq�O.�[Y(��/��-P�9W_�m�?��	욖hKq�%d�r"1�x����oY���s�%l9��t%��^&�#=�,�ݖ�:o�h?�aܷl�����@
��Cԏ:�;�k��n2���ݨ�2V+`��i?�h��Z�]��"3���a�=k�2T����h�U��rH+���oѼ�����PmQ��hOx�U���c�b��Ɔ^�h���R�ȡin_�W���v#�7�8er��e~g^�|A �n[~���)�l!!�΋�]���␈�� ��m��]�����q��C�.�ܼӺ4�ͽH��z�Z��6�F~�Rhʌ&��� ��9ZN:�R�u�[7���0��X,�}ҕ5" ����|h]���AZK�"�ϥ���y*���X^>YB��"kzZ��k��K=�dM"g��/���H�����n�Q0��AY �fT &�b��)S%�P6r���;���u����^5aC���U>�;�@�e8�?�Y�B�b\y� o�ȴ��NOA���jى����!�������Y��6o� �iR���hin9��'c���<�o%ɣumyd,�d��<�<7-�f��M���X��X��:,���i.��y�ZQ�i~���M�m+ 0�n�����h[�}e��]'SCY�����{�\�'٫2~�>�i�׷g��0������XE�:�gS"����Njt�h�8QC�u4`]���S�\Y����cl���]�^CˢfTk"�0���	��1eY��X2M�q�G�K)�g�	��C4e�QO��dW�^?�U�ՙ�j��鯋+�y'oև}�2��W�HCgC��d|�a��S�820�[g�7�� 2A/7r�ȼ=NB��'��tD��4fbiW�X�+��ss
Ij;،�`ą#��G��
]bb��A�����z���X&�����@�����on�V��cn��q����HC�<T��)g	'���T�	5DO�����%g/��޵��b)�Nwk����&Pc{;J�p|n�n�C7G2b�~���j ��'g�Mn��b-D�Z�s7�v<'aا�/ggo$t2�tÙG����0r�_�!b���M ���H�D�Rӑ��V�x��	@:�3cJ��n�mL�޴�w"��qA�>���5%T��:}��
�� ����oq}3Y;�:�iw`��@�c%"6>��\:w�}�Ԭ�����WxY݁��z&;�A[�R��h��K��p�b��%��"��g"�u�Ɔh{|�?91ֵ����������j�����dt�I?
�ݻ���Z:�>���E������B�e߼B�of�*�y��񠘴�GP���h���b�}0*mxԙ�Y9̈ݪ�6�����X��h� ���:msXsMr60���W�\/&1�K�=�~����`#��plT|�Тp8��'U������7�!�K2w��(����9���[�R�v�R�&��e<�9fQL��ѻf��/y��Ba&U'x��]cK�E�Èa���r��O����T�m���c�h@R��>�w6�����:/)�]�&�>�z��F��:G1�i�:��W�W|V�-H6h���aN�#���r#l�o�3�r�+y
wJ;V�?�f���i��&����/T������OE�^�Db�5�`���@�*|t�Om��U���(�N��G�|�!��N�ў���J�=�� Ꮘ���k�ݞ �o�K��,�>��T���j^��00M�l�E*�\;�p
Z)C��l����r��FD'�s�$(j�G�����MgM��Zr1�C�~sٽl&D����rA�{��+Y��(��0���b�=ǈ��x|؈B�ai#'��S�x��I-�j�R5Q�jj���6~�U��ϵ3��H�=�7ߖAE4�$�Ed��B��A��99׳��t������Dm����N�x_�Z�}�]��B1䄍>�p�,��-��u�Ug]��o�3�X'��YMFb�
��s����K���K����!4���BA�3� �2��;V!jDb|S��À,WT�Ē��Q���M����O���~0Ծ�-Y���M�r�n��e�!m��k��� ��q��a/�.�k[��(2���
A�#�V��̐4m���-��ȑ�s/*����l\J��eR��s���v�X�L�{�G�^��q�M���Q�k,� �ό5�Z_�x���/�}(�N�P! Վ�bϼ`����$ _N�	G~�k��)�N��b��=i򑱞i����	���^��t�Ԟ���̧*�K�3�vz&p�?&2��9<wg� ���G���b�x	�c�#h�jK9�VW����;�Y��Okg�i�#���$_�,�X�ǘ��G0,ϖ.�P�I}-�&GZg��7;B�f5�\0D�i,d�!�8s!Zw���7u~�"2~�L־��F���� �Oߕ"�O���#�sy�D��}9f0#��r������}�1�O���Ǎ[��?�8x�OY�Bds�
-�P^�ɛ�ʠ�p%�ܴ^Fぃ��7@<���M��I~�}·o�,=67u���j�� ��YU�8*��U��.���
�#�3�oi'Yl`��c����3�W�1��yiX)�����d%��X����&j�H!���-ɧ}Z�B�$��O���6�)dNR@�7=7pKo�:�v+h��l�L��O1��V]=�QT#O��<�ts��h�s`�6��t��T��m�x�x���Ʌ�� �4VX�[�[Т�����oc��|��re~�_XM�lN~���+݆�	g뚛X���A{��ÿ#_zba��V��H���)��p�v��=���M�,Fi��]uM�U ��m"�[L^��ᘻ���xԀ�gⵉd��m�i��r������׳JK�)��H��)ѫ��d��a�}(c�ug��!���j1X7�=
�s7��߭)T�.UT���EI'��<ؙJ�y�Ѽ�!�����)G�v��Ki�WA��[g5|��-l����0E�3KzB�ZPj��xX}�ƖEG&o^��I]#�qmnG7�����`D'l)��2Z�a�ѢZ�����A�II/�N�����{0�p�W��sR'�oGR�����}���Pj�T��%�l�j����N�Ft*} �4?���lhح�Q���ƶ�Q�-a�L�n>\bY��Z{����?�U��01�eg�JK��hsiq6zv|�y�[��c��Ϋ�Z�q��F/_2e�Y���B�z�� �c7J8dJP|�×�IU��6�e]���;8�W� m��Y_xm��2A)��_r���d�6-XA�)�}����N+�W��Z�T��S>�A�_��A�dX�k"�|=�o�
b���K��D��7*DCF)X���o���C���ݠ�Sn�7�B7!M葽�!�1���׳&�B��5n;f�l�&ZYU���Š��Ď�(�Z�܆��C�,�L��!X!\��ђ.|�K��s�ƍ�v��5�4T�[~ف{r��EN<��	�LnO W�{�ȭ�S��R|���o,{Rb]�#\_ֻ�E��k�[���dā��A�ƀ'��}4�������!�MZ�-l��1ɻa2�A2�3���l���x��|����ՕEa�_fmrT����x!�� >�F�@�Ij�e�7�� C�b
�.օ���ChWX8/#� �#�P��C�����pA%J`Ԩ����F���n� :1�zCI�Wz �^�Ei��+�|=��-� ��P`���;����6r�9�pLGg��+߳��k_9夣��WQ��,dg�&��BS矆)!��%u��u�=�����i��V+7Ҙ���a�Lr!�]�g�-%�Q�D;:g��/���&�?�#EU|�M���d��~��>)�#4��Y'�c�e[��
��j_YJ��]���v�R����m��o���ݠ��?�V�u���5b�_���.th���e?���D���Ab�\��N�bs:;;	�Y0��Xi?��'���X�]|�e
9S�m��� �f��x���@���̿Aݒ��M��Uj7K�O/�\f�6�Z�Q8Dꀶ;F��j�� ��A#ޣ��^z�O�h���;�|�<��b�<g�co�kCT+���H]!*aX���\H?)�{_ ��A�e#|�35a�g�_� �I��*��+z�y��J^��dсtT�1a��~Ta�M\
�a�erō�"�P�����:��7�4��0D{���SuTy-IBN�p��r���>�xF�uH�r�P���cὀ\b�Y`)c�Z�K��Q�}˜T5�>�u-�Cu�$�#�8C��yUIBbʥx�+1��QiIc��S�9X�
o_���C�?����q²�!#[;���5�����J�e�)/Y4��,ϊ�fqy�b�~%�@$�7�Ev���@�O�(����91f����:����	G<I�i��A�I�tn�	�nϿ�N)��Au������C[ֳm�!���vQÎ�@=�ҁ26͑ڹReB�Q�]TZ�3��ۇ�~C�c~a&�2�U��;�ԺE�y*�t���ɰ��/�L�Ydo�K���h����������~�!�u���z�]�:[�kV�;�#dt'��>��|�-��8�.��c'�� ��D@�i��I�Wƣ+3�K�U�֞�Y$k8��u4�vn;�6��N�G-*�YM�چ����L���6�U�W��;9f7�"��ǋ��힍B���]�<-��2�D�Cc��\��U�o���)1<�`��S�ٷFB���Q"Vn��*�l��к�����M�όL��*C��õ;��j������T�J�U!!���P�Ő�`Nv[�^r�{Z��^Ly�d���!��5����Q;]	�-5���)�n�;>n�@_үIc�7�\�������\�lGfb��`fa�&�u��Bb�o5Y�Ԕ�΁,;�<�e�O��c{^S(���4z��R�L�ِ�$�(b��%�;Ҳ����&?w�R��]�g{�gXK���u'�"�{▷x#߭��d��R�4��ѯ�>@ /������CZ�WG�\�
`������f_���u����]7{@x�£�"�mqw1h��I{O'Yѱ佰�k�>��I:./zI~8��^�сZ����0/�	����u�@8o�R�$w��8|B��U�:�Oj�e��AQD>+�&��`�I�N(,��|m3.��ܼ�2�5�)%�W2���p����@������p�2��x$���o�;������f�Ԣۧ���'�T �?�@�ʩ0hNtƨ�N�ST����vk<I(�)%[y^ss�Ĺ����AG�b�mp�=��nc]�:�"E(�&�;|N�v���;[�߈z^�uv�s��|�u��g������9����{�9p���ET$p�_ӵx�,`�N�#@i�1r����aD���pB�ϧkq�%X�r��6I�T�8X���K��૷��%R�����X��|��x��o�%P�saYq'O�ӇSUlֵ�u�r&W�
)�`6OM���%J ��V�,{p��h��43���Z,��+�����J(�S)C��_=����:�'��]2�o�AP����y4��i��L������W��Y�ZU\�(u�bBN����˓1э*+�\�+=�?([Z1�DT�v�o����i�T��b���f�q�3��Xd��h�@4�E>�b��2wD		fz�&Ȏ�a�c/�g̷݇�6��џ�x�!�Ѕ�r�V�F��5C��<�t��`@���R���	��5�
����G��b�3<UsW����\��sL;i��iVb��������5RU�GD4�s�$��dtJ\�d����[��2�{��6�I�۪��1��v���������Fk��`��4����K�h�w��X��|�/�����ly��2H�C�^}����$��
���Y� u Ό�eh&̍�+O˱��������T/z*�#��'mY:	�(0�wc�m�N� ~���w��~�T>�N��j�)����7��%<��؎�(���Kz��R���C�o�L���F9\$��#�׏sO�����u���@�e��%���#�����ҪV���M�{����,�ngrK�f���ω�h�UBhC�DrL����^]��7���F�9�l����L*�������EE�n�X��v���#�p�����5c�9as'*��<�4����譍<DRn��+�H��ք=���r�P��yK�^��ޔ\���D�弟u[^,��=�=?��'sD6|O��>ؼ�N��'˻�9"> '��%�UC��za�D������̕ch�\Y��q>բO��"�����w�FH	�a���Ѯ��o����%e"	��J��)3ލ͋�_�2��$��^aqZ�̏l!Eh0�;�y�<��|!HSu��	w⛤��;�P��6���*��`�(��d]����qY�<�,5s��'��|B��_��[Ss�Ԗ��i��\�U��8]I� :��^X=��q*�л�ޗ�3��A�&��M����Ũ���_�+���L	�3�'~!bа'���'~3N7���z�1�c��
��>�E�f
F,�d���B�$�0*��mT�8H�%��L��	-��%N"��1��x��8ۆ<��$۲u���_��ɪWd�tU��oV�[	��Z���P��U����y�*y!da�v`*��ҹ��-K���2��Zè˙8��z�%D��N#�`T�~;�s1bH���&m,C��NSU�c��ܯH�P���<���+m8;�6n0vIp*�`
�i��i���J��y2�`���������.C<�ܮ]���"t�^�?�H���S�e=�R@Y�]�Ne��i��vf�U;h�-�0iSy�K�I����s��@��  ������U�=��uV��#��'������I���ۮ���vPh���mu[�d�@R垿�S�����|?%!A[�Fr�*q/`�}9��֠��P��al�h���0��	�����qp�ŜE;��;J��y��Z�>��P��2ic��e ��L ���˴�=�Y�G,����j����Y���ן����/�4����Y�?ܺ�Č�#>m 8�鎫��BL��G�Ε��P�.��$i_����T�� !�'}^|"��B{� �H@3�7s
(�����C��]�mR�[�ԛzNl/vo����#dY"�9Ӌ�m�ժE�y	�k��i.F�'���������}==[g�OV�S�K��:mXtp�� ��pL�'�=��gU��&K"?*���ʇ1)�k���~�b`(b��FT���?.�������0�b�J���dc������(��$Q?�sP�0MOs|�
,͚�k��5�[�����D&Z������K�\G��nu�.�P̒�׸�օ�Zb���P���:���A'Αe���d�b4&{�&\ރs�ML\�~���m(�C��e���r�~$�T$f�ueH[��J�hP����z�[ꦩ��E���1 �ѳs!|�q����{�e����_��z��S���4RpV�:����'��B���I����'����޾s|N!�*��<yܷ�ܔ�G��1��� .=�Bo1��	HҸ��wpM��V�O��\�I7b.L�6�T3S��G ������«�#�g���Hl��z�ΣI�}��!xT��x�B������=����J����@�L���b�=u-�P�᭡��l�tG����'��y�nܵ� +�6a���Q�_\�Aa� �+,���f;��ڪ������H9�{���+.A˛4�*�x���|�����8�#3�!O���%/:%D��S+�駩��Z~��]���sk��ނ� �[U�ೝ��!�	[׷ :p/p�7��g}�}�{���=�T��z�D���]�A,:~[���f!�-o2a�C���B��u8W���D�n\����;1��W��FZn؎�.��+b7hglŦ��ą��T�d�S�S�G�_:*6c7���(��7JOL�ϑ�\qrC�L��6��g
i��h��3��x���w4Ku��(��M8,�i��TD���m��^�;X(l���8�̼.2�H v�t��N)О�~c8$�Q�è�{�]a�\�н��NɎڂ��$�X��T�ﮢ��s]�Du>ݡ�}]���J���d@9� DR�_{ߛC��u�J�����£a�&f��#Ww4)G��}�3�p�xT�	yb~�(��s����\�$=��Q��y	|Ss�������e�c����m�{@zT��6�����z� �Nd�,d<�vn�՚�e0[�����9?���,0��,Y��^ZU||�c�$,f�_l�����04X�!�E~��Xx����phuE�|M6�E y��Q��V~���ᚖ��\R�m5�aƥ��3�AaOJ�L]���Qe��>X�$ `%�p `R5�9NÆ-�ϸy+�?^��Rq@�]�ǭ3����(`ٌ�#���ՁΕ�? d$�Ǐ�o`�ٕ���A�Jļ69�L��\dpmeO��=�̚Q�����Ya��R�ҦЉ�˘��q�L�����8��NF=�=V�\����m�w�Ҽ��sUN:��c��H�sٳ��q�v�j����8��,�OA�SK���Ty`�΂%?|����z�'ɚ(禗�VPY,�-�*R�B�( 5��O�g��w]��B5�<k�,"C@�m�SXS�gP�����ǚ�!��������\���a�A�!	A�SdR�����8�Vd�KƆ�g��6����Z*�l#�R�i����&�tk�v��t����i���وD�jJz-���/�N?�(;��f�qA:Y��^`u0	 p��}7�||�1h�?��s�	n�|ञ2�B �o�bE%7#O�t�$� =������+�����<���1)䇅�U�J�!��9�t�
_�_�N�K�33 ���h;ʖ�W�_��W��ߑ��&A˳�5=����Q�k,ۇ ���c�\&.(�5�$�&�eU<�'ß�����K�+	$%��>m�`�6�O	��䑺���J��P�Ȅ�x
�Xx���z��x;hv'���O�ʾJ�)��Жj�D�"�@S`����!/C��p���I�AcQ$�Eji�x��"�a+:�]E�L #���*є��A��\^:(z�;�J:b�c^�𹙰�r?�zt��O�o�m���4�*XF���y��� ����в�uC8V)��B��
�F"N-hyRs��upX�W1YG��qT�k4��RXI��~��XM���@ψ��z�NEΈ)�y�I��֣D��Ů@m]�N4��f���D+���z����I־�a�!���/]q:+k]��
tl�.;����g���p��&�y.�7�E�|���m�>Q4P�ǦX��?�7�m����3H���-)�ȍxd���o�m?
��r�q�!,h>y��FP"��� ����������o���N��d︻w����8�P�����Ů�	�ÄH�V@����'yxf���Z�d�4��4���E&?n��ӕn�MO�t��H�|���wf�7ڋ�2�ݵ]B���K�r.�-���K"|�e�@(���B�P5�$�9�������VȪ �v^���o�U�XRcT�� b�2	X����+\������W^3�pߴK ֛91aI������i���\��Q��weF�d�t:g�S�%g�dΣ�3���o����G��S��#��^N������,�b���9�a&'4c0��w��"=���,��ëQC�)�&K���z���5�B��Q��!����w�&zT�ض"�z�Z#)�X��@C&��S�3M�r !o�����'��U!��[��&&I2@��7��dD���uu���	��%5�WB�?�����'X��;8D��3FzB����AoC�^X��)��"��5J3��Rq+��2g���&l��i%tbl�Yx�'�.��X�����xVXk��g�k�0m���(ǅ	ω�㒣޶���7����/;!��~G����T2�)�4uT��
Adϓʏ�kV,�p1t+����41�gy�X�������Y���,L������8��$Ӆ�Gӓ�oY�X�(!5�]e�?ݐOfQ����%z.��P�\�<rn�u���@���/7΋�KXr�P�Ϛ�l��U�T5�
s���k-�$=+����ӻ�g��70�ٰej�;�$1�Jt����TL�P0��k����)'�h0{exy�V�v�k���P��j��38�u��6|�p������9���u��#=�Hi�`�鷠jX�-�#&K)|L��H�)��~�U���5q��7��Z㏧bX�|����]����Iv � `;�暁{i���Azqu�~�i��?5��l���6�Z�IuBcg��F��L���+U-A�0���^�;�_Y�Y¼Rpg\r�7�p����G���b��H���A{�ʚUKN��7� C;|Ё(O�[�;�)۾�9��,����K�[��y��\k�w�9?��L�����ט�I;]%��.��R�K4�� �(�0�Z���AL���(������W|�V0/�Bq���8X�n�Wȏ��>���N̛���k՗`;B�0�(��Ű�� F���� ͣ��-�#g�Q�5�B�0-{a~�S�#�A����C4���R��:Q}�^ɥ���u��D�ch��/����(ʫ�����|�8,d�Ҡ)��N|Ţ`��.	@���o�c�>����%�\O�p�]�v.1��GN>q�ЭU�<�b�~��Ȥ�)tgS�)�K�~?Cr��;+R6qf4���]M]~EӞ���:n�4�����8��s*K~d��Uh!Tr9t2w����;%�+;�o�>�})���!"��Z�%2��\n�5P�O��n��r77��b~��CQ0� ��R���r�?H��v�4�� 6���0.�>�Q��yGq3�ݮ�_0M�w~%�&EV��.�B�4-��G�`��`��'�-w�����qMc|�o�?��Tp���v�.q8���R�]���O�Q��������Q�CHd'1�,T8~h�*��U̫X�%��M���V�ɷ������qù�vk$�:#�?%8q����҆�l}S��>�y;#?���g�2�x+a�Df������`��*j���ͭC��o:)�~�$�kWs��	ё��R��霟���d]��|T� ��9;�|����^�c�ʑ�V��Х.��ǎv-�C��� >v]�?;�A�{JK(r�}�3�� -�8<.X~S.�b���9��s1<�t#ɟ��%7h��2.�Àj�-*-G� o��}й�K��*��ɼ�V=۞�XJ�~�C�O�uD�i��A��B�ǂ�䦈�#�!�*�H�AZ�S���w��j`��m^�A�B�A`��~T���9e�y2珺���|�}����L�^Aq�ɣ!�K�G�i���c�՜����)�^]|�+�P�}�S�[긼:<e��Zl�ށc��i���0�\��m�$���|Ǣ��ӒK�(hQj�[v�����3��4=_�Ѝ%�i2��(��}�zw����aF���V�/A�*�&�#m��:����x�dm	vt���^��<���I��|m({�]����5���/��a!5�Dq��t
��[�w6�>
��M,s�~p��O�w����{_D��5�۽������}�����ZƘ���s��g��C�l��A��F�d.�#����X���>�܋)�^.��uN^]�̮��I����L�	�*��5�Ų.�vS#������'�����ֽ�wm��U1���r�h�(sU�[�T��'�N9˪���z�D�T���˪���n�訑4�=NndO��C(U�֧x+�hj�YFa����룍�1�E%$�����͘����xH�q���"Π$�%jdέ)� ��
�~�S�9�e&ZJW��[q��)�_��`�6��+���l�E�>���V����M?��s8���2E��´dT�5�q��m�9==o��h;����n\����Cg�j�z��?�cRR��4���1��+v�4i����R+�t�s��Q��F�|�	�[ς����L?���ڕQ�7��%�[���ԇ���a��-,����/F\�.A7�B�r7���vD����N��*0��Sf��?"i�j�&�'k<M��nY�Shr�/���SBl�+/�7�4͈��jr��v���y�z���"7���P�=da֔�?�wB.J	
gX�fH�]%�U�F��K옼l���j�,D�!"����G��������-|a2G�f�����5�j��� ��[�m�I�RgT�
��
�:�
p����v	J��	w�S����r�~]�'����汏K�2�<Q!k.k��	V�_��+|���9-�o[�!�-�_��A��2د�܄h#jȞ"��}j	q�쵹'��V\�"�.'0O�E�d-L�T���Fl�0XRr]+%���O�3��g(�a��I�>�<�1��]^sx�ՙ�=Q�3�����pW�J_��jC�ïr���iێnr;M�R�m��W�W���0�Iđ�%h$p�d7����sMd�a-�ۏR3��,���*������W��� L�$�	��"����^�L�R�Я�����Vfb����:&v���8)^�k���Z��.�5����{xTjq�����p��/�{O{��p�ͨ������GTw�/�_|��8q.�37ĝ�"#O��_���!Dw�l�{m�^�8j�R�i�=�کw�{gL�6���C4AE���a�I�Y����Bs��Bx��+;c��&w�.S��0��Me?���bꤔ���y���T����y�(�f�f��L�&� �-��?�/��`52�[O��� 2,2��H��Y�Ю�2� ��8^��v?�:�=6387b�I@�D\�b�0K�t��\�Z;İȢ1�wӢW�[��n�Ή�8�H��H�9-ő�	a����u#{_5��l�(l]��dp�����ET΍ֳ�D�f#���c�w������s�1��F/œ�m�����	������}��#	,�彂�*���9`/���	$���\!��&����7�If�'���ȻF.T��m���a�q�Y��:1z���T�ܘ"����N e+<=�9��T��y�`�n�/�D34W�ϟ�v����[뉞�r�|��s{%Ӄs�{��O�J����#���� �7� IK�PT����F a���Ze�\�&�Ǧ#����9[+�0��|����ا��E���2ج�BSd���_g[�,��MT�t�Ѱ�e}��܋It�]v���!��B�-̠��;���J1ȴQ@�F���@�d�DOD$󛑃Nc@���b�ni�_�L��3h�a��+��M�פ_������qAé�V�I�XdB
?���\_� �ac�|@bYk?RD�`e���^�"��jK�ˑW��FU�Nru�u�}�k�;�˨5���+�O7=���"��A�����.���0ϗ}l��mo.9�		�4�zRl����)mTׅ����0��uŇVJJD7BI[��c�u�%Ϸ߁�8��!^���k�4ƶ@-W�+!�E&�@p��ZԦ��
8 �n�4I��ϳ/`Q�{5��c��Ic]���(p��b�I�3�*ܮܡPZ>���^���k�q�-7�b����><{x�j�Y{�X�ڋ�*�����|���b�1��`W�ɗ���:��X�ɶ@4�ۘw�#�'%ɶH�Л�o�Xi�u�ـ���݌m�,`�Ԛ�WE�%K��(�A�"�cz�V��3�Y@O���f���G	1�v&�,5D�8�jcY;N�WY�0�\�,��(̋��^���N��u��`��xR򎍮��s+��$�۝�Z��$)V;JJc���[`6�,�j��0̶�`����\�0��ƢV�	�x��ŇX�8WFV5�c�d5b�qW�C�n>�Ţ/~����xBVW���[�7���[�$t��š�*�*#������44vfͦ���2��t4�2��?�x�:���q������L�;��i�]�� ��"�l�a�JJ!��\�2��b��T���1�A����)M�z�-�r�������uC��|��n��=�G�8�b�=�eh�lh��Xx�mҲgI�~.Tp0e��Pʙ[�'D0��P�]��)��B��<Ɠ������� P��Gt*���$�0�%/w���'O��۔[Ù�!-�?��j�Ā��;f�V��$�F��> =��c�����/8	w�^�O�o�> ?2�j������^������@�x�نcA"0�t���k�Ȧ��d;�3��V���c�����c�]�I�W���QD0��<k[B�<ٛa�k�M�*��h� �6���5X<�Od�(d�زeb�gx��~�~j��0���M'dyy���r8��-̉-c�2g��qL���
����O���U=a���nT�J'񮱰x�š����P�$l�z��gx%\5Y�E�FT� B��VnE~Va��Y����Y-gc�_	����$6�%�OH�����n}����8�ǔY]JC,G7�K��4>����ZKU�]�x��#��lU`Z���ۻ0�?+k�w��[L�2͋ߴ��wvN>��8F�7����,�ou�AC̍'�nJ�L�3Jd�������Z�������m�H&{��J>��̜�[���E�{	PLN�u�!�\+*����CT��ڡl�%)�����@�[�� '�bˋ�>��i#Ŗd��,J�#�5e��/�������S��$�+������(�P1��#����\��Z�J-#o����ݐB6)����� ��U	o���4N�=�U��:�})���u�s���'E��8)���Sݳ6�|���\j�6��#�RO�~
�V�/��Ƀ<!	�Y�N�l��X&���}YU�V]����AJ��b�[(���)r��]*��d�]��{�q�C�-��Ud�c�O�-�����K�6y������"�l�"?�DLn�!.�T}�nb�����
sl�:�S{�n�P��)9�N�p5O��)��lQ��$�vwN[(������ы��Q1��-s��!_��\/J����tB;����S�����5�����>���h�W���>v|�[s��D�vs���8.��+��d=e��Sd�(f4��M�ޭ��6��4F��"N�4;�yAZ)��4u+I?(���ck�̞��h��YH�Q��E��*���U�<n����=�����}��ގZ\j���7�FUh��k��nuf�������
��t��g�G�Š~8�S��Q���[>&�M��lv��S=y��<4y[�<�H�N���4�{�&��-9��1�L"`T��:]w!�.*�4 �d]�瑚��e�j~�����#����V֓��B��UDs��_�^Uk٤��[n�x��QF=*XX%��ff��AI=s'�OX�t�>��:�ዿɡ�� �l������I���gny��3�Q,8���w�����eJ`l8V[�y�Dו�,���N fO������,�������gn��ןrP�y*Y/դ�xj�et ZL��1�v���¿��^�qG�';��˘%O�DGV;�8&D X�B�߷=�^:�qlR��vR+j���n�V�r$��)hHV�m�D��P�#��YY���F�"��L��EZ�u�� ����f1�K#tf�&�xP�o�G���*�"�j�֨�c� ��D��o�]�l�c���v�/ Ɩ������.|���f���	V�}\�	m*�	�p v�(8 ����+W�_?�UύC�KGm��ХM�5-�/&%��,ΐJrз�3����`��Gf������k���no	p'�m����i���G����0m?���[F"�����Ψ��$��4|7(��+���`��<*
|�Ri�0�5G���yb��7\�p�D��iR
�k3��03u���j5��-���@�2-lf+�zlݩZ���$�~_ei��0晙=��ŭ��FA�N���H�%��b���@�0��z��P�%;<7������Zl�l������o�̴Re�\	���S�3�]N���5o[M�}9�5� 0[R�<|ŲL�����c���ν�e˗P��+�LwźO������ה�g�>��.���+��
HZ��	 ̟nE��R��1`��דKg���N�E	�AU��nW;�l^���Ԇ����MsTt6�/V1��:�����F�M#&R���9$ռ����y]az��&�/�4�Ĭ-6���d�����#ُ��i��"�����%9^�(�ʗvJX�J�2^��7�,K�?l�P��	~<�0�T��Ʌ_L��`�b{q��gjO���.>��q%�����u��w���(rP�
0����@/v7%}�H�,j���Ǎ����SFP�7�=��^�M�R'�!��2a�x�SH~ֽ�NfH>��v�JĄ�P�ٱ�{z��3�p�w����6a�w-��y��F^S��� ��myGX{֬x��6�qJ]ѐY:����G���L�=�׍���o��F�m%��~Z�nK�=�<�$��A�9�Cn^�HւSB�?��4N��F~v�]]$�ۣ8���􁉞���0}�7{����Q�i�F�O2Զ{\����@�ޜnAD'�g�ELJ�ThC�=_R�ew�76����	&�����)^�oy��¸�ŷ��p��T]��=��.����k��3? �dsBO��*t�Ѽ�:��#4�$�(X�/�E%���IYޛ�T|t%j�w0�`a��d�G�NJ>ɣ���UEݢ��c#�9���u���H�W;��V�FFt�8����n�T鈨t��X��@��UI#Ɨ�P��Q�~~��z�&�K�wڃi��s��rD�Y�m_��0H����q����V|a����]#�M��	���6��x��p��eC���Ӷ���*�>�a���˕��z~%|�A��*�k�҉}�{�(�YD�n��;jX�jͪ�Z��ܞ���&�p~�.]�z]��[��טjUo��qݢ��٧M�w:'s��/��S��k{�z�U�H�L����n�w���W&�q�gG�,��>�Kp=F����W�$��=�6i(8�WP�yc��	�H�Z���r 0���*�w�g�W�����.j6��6����{D�(�d��&���Nnlh�j�����F¼�6��W�؎�D�v����@,���i�����y�e��w	\�qO$d��k���>�Y��*�șY��|���.�>ˡ�M,?�Zpķ���w��x��a�=� e�7��Z~:Ig���")��qtܝ�]RkY��k�����YE`��9GpS�ҿs�I�Tq3�юd/(b>�&�=bG^����*��������k?�
�C�}�+a_�e��n�$*�4�6*`�?.�q��}����ϵ�\��O��#��	�z/��])�@�|�����'k. ��k��]����Ӯ���t�X��LްmU�1�>ŷ��6Yf�4C��{�f/p�Oi㇙���{�@�AH�"��O�Nმg�kg�\�Nl%m�w�J�`�Z8�k�1M�
����V,��̄����}����=ϥ3�����������1
v,+�?�X꿖�fE��u�:�Lѯ(��-l:��Y�X}k��( P��*���S���bU��&�¨�jt���H��z�萢$��R�mk�Zˁi(�D�'E��p�ᱡ�WÙ���B�CcA��{�z�{��vkT<�,G�7�@A�x�_4���zሒ�+��{#~%+��P�1������i:P4�b����C�0��g��ʸ�:8��|X���P�h@�F9�	�ά���#�?���{�����(P��>\��u.�-˕���܁�U���7�4"Y�r��Kl/g3Bj�N�uA�C�nt��{�H,�&'�X��z0���,j'(��P���1~2b8`��(D��`��+;�۹����*��H�,>qU�P��ؽ��[Y.lt�z��8�l}���}r�\�@�Ѫd��E���R��K��&��O�2��ǅ�hU�{��2�6�Ȳ����>D�)B_�0n�� 8`K�>	֫�6q�=0y�Z�j^�	�^������ЍXY�tG��G�Ev1b^C�!�n��ԆZ�R;� ^�Z{�����͸IV`_b��z]-J���Y}5�s���#��ޔk��	��FP�0���|�_��X�U�ث�(P��<��N��T�E�\+��um��r]f����L���{%���.Oޔ��o��3����o�0
б[G�c��Q�v۫��0�^..2�XYn���t��H2W���l3U��>�
q�
��v��y��F��3v5y� �!�ۍO�F�hh@Z�\�PCY��`�f�9���T���v
�R�>X��d�(���;cu�5���S���z %�<=�ݼ��X��$�5������bA	�T���)�p4�������ܦs�r	!����i�V�d�v��ᠰ*��*�Й	_���K���~�e�}�d(V'���<�j/c�i" n��3��N��h��%UdXk�H�~�>�N�g{�n
7� ��;NT�]�h`>���D��>��*s$6��z:Acb���+�;9�3W"��)�<)�i5J�O��
�l�D�!�
��T'��s����N
�I�3�����m��3#�_�v���ݼ&l;9E��'E���7���F�#����Q�ܶ�V�Ǎ���q�M����?Y�����Ț��yc��_�I�۾׹m��k2q��F���LK�rF�Kƨgbү�u',��wW������x��,��4��p��e_΂��{�|�㝾�_0ވ̤�	ۡ-���g+9���w2��{}
SIŨ:�Js�;�Fz�=�U�sf`W��Y=��0�φ]��,�@���,g�^�P����������Ts�����W���K�`S묐}���j�m#���7 �LY�cS\��H[_O��c/Q{!�1�o7�����ȦC �6���iBx�g�^�?NƩ�Vr1;��{#���1�����w�=�?g`�lj������͎r�p�>��������:�ٻ�a*	��f�3�{>Knkqo��M=`e�A˅�>C"}���f����y�xUxpCK7=�|�j/i��$;��4.I��x������/y�[�����mNq�*#�w�/���9Ɂe�{}�s���;��I)��\#�I�XRΤ�Z��������=���3�&�K�Gh����~M �����5p;�Ͽ�H��N�<'+�I�uz�q�_�)]��U'�a!7@�p� ���8f��M��{)!�A�ui`�D�(��m�Ol�91�J$Ѕ��y�c髗X��������|�
�0�E9˽�[�^g���r{e�P`2ڈ/|M,瞣�����(��y�辷l ��nΤC!���r�츇�.�i��-��