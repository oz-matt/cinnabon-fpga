-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
M7imKIK0cSbxHvAK5mElQtZb0XpBIwwDDyk2hlIiPFahkQAWqLhT4G5LGj6+kK2VEpecWwEPXxoe
okpqgDmO4LR70vs+GflaEbOllfov8UFBmMvw3dr7hNUBdh3PbAdeOlVQCtAcnoZtk76HLcakZbHx
o2KofS4gYSRAv85HfWxuMK7tSMC4wjWEby5NdkykWVVZwlD4377gZ0CjYPuUlCrhUIKv9uEpmvNr
YQJ/iOpVzFfH0xeUUyjsBl72yIr+5Cz/NK6jhh69cR27I1gZUat1nhBtIHR+/dKPvKNzxAfRaYth
uySDAFEDjb1D0kCmdGjbMx2KMDrJogfDbKg1fA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 5376)
`protect data_block
MWP+Ex1dPEzrptD/GhGMMqSumhATkR+o99jy8Tv9JJIUfrMlVXJnvshxJRmidoXLDJJYFuNRevOw
uUBpj6C55b8fxrpz3VXMUrVKJiKTx62/MxCbshnSGfTMuH7xOrfbTOwbOXawuXsCAxFVyRqLmSnA
K8I+Wna8vh4p+th5odrctpmnY1cNwYNMx2EwE4+KWy4NX0rUAvdc8FBJFZd9eg7NsNOSAKaKRdfb
W4TIrrb8fVgUOawzOW0r97HfbJMqsUmJyK8JTBUXKk/NNoO5Vh0SSZ6maO/kEz+7eLZuSAA+tMGL
0xKyXs7K7xUHBKisdvs9nDXLi90YXUVLptYu5bm4qdYmd0lerZ9EDr0PD7pcPgesTrM7hTPw809R
0swWz0n2vYRZtxInj24FwoTwNSmHkxHIznB78Gjj888qjUkfrf7hnnxuKIn3kst4G3i1aZNAbAJs
bCxTyodPbKP0XCV02VYJMbo/5aoqp8qPEPdsNFz2Gbh5Dm79hy8I4TYuNHwtWo2DNlLfqwmaNfIr
T8dK+8Q5D2dQlwUfeZBXbuwzuFe1Rj2ytJBUIt9TnzA+NSAwGQ067EA0G2MAfP4XFp2JH0CRMm+4
c6XhdtckOYpT36ISDqPZHOgUwD2n7IbiaQQNF7Pyb4FIGfCX1eGUe+iL/+IcC5pue92/WLpogzz7
Bcl6Xc1NOKhOXZ9HjBgRHjJpxiXeQzrjPx9v/M/UQ4emElrUpH/MHSOoTV34FILgJivmI2sJfUUA
q3CSSJTaixPkp3o42Cbzs0BfpAyqMMb+PDmq8djo+0YJqRLOFrRgd4RIX0K5QI+mIPYvB1YiJWNr
wCHxqhQdpl4KMcxMkqwj7qZV2K/2m/kaxXI6gaSFqynO/NCy+Yk1ZNGaAJFle1Xy+by/2ZMUos+f
Cfn6C/ALgbzPxrvvGbsMh1dhOW8nSD0ASLPOhdM4/IHURu36wJK7weRjbia3k4nMTgjjLH0FqmjO
GxvlY3lyuGHfGdM8x97T8ANlsoC9fcmznEGummdPvHTjZv1qFkACfcx8/PeZ9VMOjbgWwa2PRz7i
ob3cKs/ofoZm0Ykc8bOPLyNPGy9zB9Mpj5r8OOTw2EWmiC+BKyJxfKoxrzxKj543cEJ/X1eF3Mmn
i/20xwZpUHUVQ0VnwcWuVGt+CA6EC2Tgivp5xq/7rCoPzxtFYcYpvbvQ58BfAXZ7Hi6rsabe8T/y
G8YJjYzXabZ309l3VOlN7rWrM8IJp8tbcLhckrEC4fDxBg8rRLus3BHQeonpLZ7wWb8YjB1HQ2UR
EHtjZPhXghVfOo9QefL36sWvPV7XuZVWX1dFWt90JIUdh+j+wBI6/uXply5jZOaGo1JBcVqeEJmS
oAYSbC0AM6g8pn4vcW7U/eZLpfdyAWZvddtiFTiLmzLGEow1X6OrOKhF6+zuSFR06W8iBmX1TOKE
8Cg/N1QfOL6rdBWRyfxdRUVj1GblF4LfB4UzQKLB+pxTxJYMVDWg5hrSmGI0NOyJkMW2lSirZ1MX
ytoppf9HtghaixDc7seTWdvEe+rDRuhT4OryBj5gMXiJulMe0/hiEEoZ7bumHBzPBakbDhGslVdH
yRvFZ9bZTCmiptn7WGDx/1RwWqWNAc+mTFDQOFbZFj6Nlq4hmmms2fxhqwW9ZkRoSgdeGyOzzfFA
UMcqv/6pU6UB7cyGKM22FzGKAKx2/u3tBFj3I049XJkB7EKzjmreNYvXH7fzIu6cxe5JlGGK2cH2
xQSpNHz+MelIYPUrzCplR+G9omMT6pNlRYY0tW/fkipout/ppyU+dkMpXxpRKFonn6XP9egsORuT
99d/OqZOYyzMYVNsaLAF4psUdW24soqgAm3zmiJmCQvej6P58pB/EoOxXMDwt4vCQ60MIEczKj3n
BrlYKEnHRUoJ3ttuHhXTvREzk59+56PaOcBv3s2qdvvgsFFf7TlmCl9qtaPFNQkPHCpLQJbESV5+
Sy7DraQpN4p2yx8GQm5cEZqZjlCGV/C+R2ScB183Y5vmfAz/bor0CslEEStAPmSRATQBNIHetRF5
bnb6T1PefnMZ2rVlQlGjtLz/Bq+7G3HlBB09L7SW9JI3xUa4U0c46KYQI7v62donH6eF64g13Tbs
wJyYGUOIyzHkJ6Qe3RkLCYMkEJiMzdthz6fq5ijJ4cLnwy+hA0J/AwZwUzbjbqmHsDNb+kTef7Ed
cS/FFdv2qeUZlnoyt4I+mZeuKkj43Li3ih97BKHpvM9CZl3l28STiF6Umz/M2LEAGWDIe3AFGKtn
OQPanYzGqb0fgwEsreNkDnpqXbhJ3Ln+4ZlAVmobn8LSP0aKRwIs7LusLecBcjYrRN9ei1Lu0elH
uHq2G7SPVaIKMcQQzvmJe8EsgJtoTinARMWEaW6JZdhpJHs/hlTbOppAar1lJoxvF5fkKml1s5do
P1XfoMv+aTxz/VBfeYH2hE5wLZudjw5Fl0NCBJ4pThgNasvwA2UN02dPDJasOHRWXeKXSEIH02WG
s9uueyTrqahf5VHL3w/M0POa0K7HOCam7FmADNqt1cR3FLQqCRKEaF+T5lA01ds+xLKCQAsR6Fzi
oS9DkIk98mkqYzC56bNTfLOjbIo6wq/tDF0vuVdYhA9FjgA6w57OkonErxylcD7gB7ROEnxB4/1v
ltVlT8PvrvMRsyAlaL9xMSB/1rIQ1V+rYwBLCE07bdWW8zQxdeuSoxXxw7cHvSKHA3qtqjba04U3
JOipJh/ujE61s2RrnhyR9WFi4U44C5vmHuXxUvnsirGpLG1Y00mgtgfnj8w8IeeRot7JDBTfqCAc
N0JVQcwMq/ydRur5TZ9HgYU9KMRv3gKHo8MJL16pNTcWt6wt2D9fITwMbLTgg2QgjNyHtAmb8Agw
e7yBJORjEfy2ELHVK/vhiXi7sbpc4X+LyLRJDa8i3D0+wAG0kZjzHjr1YoVfIE4BlTm0VZockNTC
cEzqMrZAK5z5mfd4p3LyjmuvVowOzgtsEn4IFgQsSmztEnezifsxcp/31yS+ijIg1eSaJ/8G4Vdo
pKRIGmLDT6dH0GWmL/ZsfPP6PEMu6ZZRvnY8Rn0hldEjdJhDx4EsFcvluDQa9Ubg74agAUabj/N7
wqvRgl7t6I3zCL99bwmGJxpfSFd/HN7Nvk5Q0Oqfr3PnINbU3ekGaMieQWt+n8PHm0ug2dzRCvfx
U1R2AcXq2o1fLoEoAWmagvAk02Sh8fTUoZoVHMBodvsz1MCftxsz00OuByQwx6azdN0gfb2S4rZp
bkx5kAChq4DvYyDucn3nrZo8m6vd88Rdff5EJPzkIAtg4vubaytXh209oJm89800kLOaLpMQ3TzG
wsAG0jsQZTa116UXq1ULAP2vx0yKbIisCDTPeEXUX0gNGV+TCCX1uFZtXXxYDFFEYd72l3GKieVe
sl7KKjw8pCqx1WaMEvfy+EiD0QpG5i1Kn6CG7GwcMIJ8tTcE1EYMNrefJ1+evDtEqJ0fGZOlI0Pm
VBnZPKcgP7wv6KkajwzadHFecACwnsMbFaLNvTwcGd4jZfPSXh/cHBy9OSjid4JV/Ld9eOW4kQo8
AckyQ5oLjlSQ7OcvU7Ck2ETxvyVe+8E8HCj310+yZiLHybZ2O7+TxUymhHnqQUXLx0YoKUjSxRra
vJRSA742oWNFdiuHYJpTj5bDJJrtFRsPUSoPwmTfS8hErTbB3E9Tl/stuUhKJz18t1wSMRMuDbQw
CjhowVwY94GAn90EacLXzTftb2oFNKDUfYjbzcMzfdfu5L9a4AdXfcHZeNFadqzcG0oIgyVB/FKk
QPm6sRV92cB7kBtl8fs095mU1Gu2dO5jWPuepcWtxZcZzB4rVIkOyuP3cXXEcFKEfp+f35gNm9gL
F+2QdkR8+sYZeoa0DdiKzYv89BqZh2FxcbJHsP88LpkiI9yFHTCP2eZG7ajdjn1PMeMenlHgqgAA
KCnc8UYfOEDdtOieBlXrSMoa5b9xwtwWb5VYP+W2RpmpNYHF3+2k4vU7sCGcJ02VGQHg+tFs3iCQ
Xr/yrsqc40NQuJB2e9BAsxouRG27Xze6Two8RZTA+fSBbxRTv9WJqWUwRMxjF37UpigXea5jHmVc
AIFKPJV+dgk8u/6JxNFXfaW9m6NjMzz3d+/S9cfId0kSWxB+/DsGyK7wp48dJWFoOIbEyRR7yBiS
mzmEE3UN6hjwFqzmbJxrJCyMpwRILLqc/FT+FJx9z9t17cNlhn3Ec9hL2JUKe1/mPWnFc8pdET9f
/FYvWffrzfQGPDL+ZmRvonRQSRs2H7R8Y32ADZdfSzPaqCxht1wm7aZkw5APZfqAajheg4dYZiPl
QRxQkZhKsZeOY9CTDpkn1XXAogTGaRML0quguTnf14guI7KgjhYZ+W7O5NLgINdcY41dFPl3cZnN
q7QvFcBUqbTE/KxjAt93tWpF8LdV0a0ooSZcvKdsUr5cUr2IXOhn/MjqymYxLvEL+SpuJCf8TtB9
g+F7Bl1sd06nw5af7tYTnoYJyw80TLAYvpKFVrYj/fGghS3z0H3hP57t4AEM5S2INWKQ6wBQ2g7b
TyerA6toKR2WumKDw4oKbtPGzMf5PO+K9TBVRPPAAVNY5RmKWfMkGi7rT583nK8z8i2ykntxIX+3
iKOkd37XpOFp/Q0gJlYX6jPeDuUMej8BzVAwWo2qmjgjp8y73AFvOCRTUeKrxfUUqd0LUFPh6PpM
WbGZtdHq2bmiYuPsOLfcUBvguoIdNxhbwAO/DUCg6tCQ3x2i2ST/fElsNwx5VAZxXwXluulaqPzz
Uf9TO2GVrbxCHXuHLmcTXVccApT/W/ss2jX/I7krOz647srF/CJ2kiWNGuFVnf10ekFV0W9Q6P6Y
P1Df4X9qvQDpRfrdx/qQo/89OS8CcAsKl1VCiJFmpQrytJK7cpjwN7RC7uuE8J78BUc2xtTDv987
wEXPo+ley1lMk7uNrg5QK1SkhiNW8P22oxp6m0ZMtgtjID7CO1NlCQxiVTJQeBgB3bvxSsy52YlR
mt5n9fOg9U+NVtAZNiTREraTv1GjButZg6QlXjN1J6N1T6fPkqPaEnPIcAAvioDAU3A30c0H0y4+
sEosOgdSTlsns5IVWqL7RJVhtPQ+//OeiZQg+ajyRd14lF0PL8yQrTO3yU8mLv/ky4XVzWJ4q03P
wRKXunDHrk/1L2ovXTGzELp3baFNEC3x19tv68//OycL0/xCmBV39uJSd1gHY5yCQXrSnIT7rB/V
xm7aRyqkDCHZTVgT/AHyBhze1IubVf03EDzFIX+zAnUDZFGzWWqeTAxewaZjtr4TO/jYmVQ6cQfU
KDiSo/i3Sz08VLcPIe9F6TS7Exz1/xyDTeE0Kzf2T1chmCimNCeTe2oQ71Go1OMoOq+xKnZ6Xl+e
DQfXISCr9OYCf9f7Kt+Ox4EW85JZ4hmBBaBISSx899KcL0LG4DcO/F/dmWJf8yUO0afxBdUJr+rm
R3xJqqn4y01/W/Cx3r9cu/lPRUX/TBNKhGfPW31zRTMGJ+ogmWMjl2Q8xVoudFvnTQc3B1HISxbG
CunKGmULa4YQh3pyjXtYiXXhH+As/kHrQjMaOMg9yy0/d0S4UYfnY6Gl3mqhHj9oXfgiwPQQABAj
8gDxw0+D454hFDgrtf+qydHveAMNG1LbVpeuzfUk2wGyGje4ANGdN0qlFTZxAqA6bcOuSSaWTuV3
A8D+DH04m51AKf15nDBgUQ49nfFN6PiuyaTHdWhKgQiuCC4t7aKhUL1/gFIxJ3wO0jqQRYBAn/pc
gOUDmLhPqgUgi2Q3rgRxzvx30F7n2cTEyyws3zZFVOJLgtjDjLGqKy0OqYbdRRUjlzuzt7zD2pJz
ZRZsNwkaXdpSLx108Hfa3SVImkyjxyZA8JoLqzcbZsYZWB0ZakbO3HO/re4TidNeFBaRntFLCz34
JXCyuPwsZJQ21Aj/T1fE3P7ejZbEsTiIWa2RE6VR25jmsPCViT7vZ8vn/64WT9Kbz/INUKYrg6NY
DjnG/c0/aZ0iMi99JH0MoFT+6lSnOIuCxlcia883h89bn8J+IDK2+RUv8Xk6elwMxWTcHMYBAVlG
LNFGcX/YiM+y+iEAFpaVc1mfKvIvZj6xUWKD13JI8S+ujDXWE/phTmaS4KJfzhXsEpX+ncX0URbq
hNN/9t+gQRczA6nt4WkaFZf7UsEIasrc01LaeZsEPD8LNPHQxPeNMITj9k9Md56Gemk+TXkfotDo
YyDASxGQk7V1WQ4sb/EjJ9tC/UDx/F5+or7Krul9Ab0ij4swPmvEpBRMTLpuomExjXD0shOHfFxs
f+oJE5wITsU1baHNJn6oEfINSGWXFm+XPY2g/gkKV0p9dieqW/N4T/KmYA+NGYUdPLb6Z+j+iXiV
FZKDD/HiHRBTdPdxtc9L0NNDCSi0BZy8E+M8wm1x3cX9bHP5GJSQUbgWTaNJuAHfqsZ76QzdIMQY
LFzBpYXLeKOquO5dpx5lFcETpRU6mxQ7Tgt7+y4AuMVmEwxXkjnlAhWhOqHSAogpCY16kZ02pWO6
K9b3QIWUIBbeKS/9YvLo/P6SO7asMcq8D+AzaC3OmNp4PMg5FbKQBv5zsz+RhLmeBNR5o4d25wK1
Qr3f4OGxvh5XicP2VZJ7yPrjaEaUiFKkq3uWMUmOrDriZq91yDCfZ8hvCJupxNaVM+Ld1jr4zsoj
VhLWgrChTyn5eJVa1zL0zmVIJRifbri4tcAnUf0pbk5rYJuGiAHoVHJU22CMg3yaL9CM3eGiz4ip
AuC/UHKfo3JunXXUxAW79WxkrJ1JLXPJeZhJd4viFuHpXvO9LqSskHVqRR4g5qOLieE4vBs9uW4R
WtSXNCeqVWeoM1G9rhY1kL0iSsHnqvZr8ECAKxRl3iPuOOin/nLQyATBSVV9L8paghC32MX+HMs/
wx8ZCIHmVICtnzmnIu1myoWbkJFZb+QpdIKT0tNxweneuvu763ExR3RLOSgXhhQgjcyyhtKNEFWn
NWGy8PrJLV0QAzCaTVgxQYgYhuYL9awJDjtC4LMxYEfeABN5AU68RfKEwfFT+5ri7CG7nPR+96Tu
GL3nB81wXFxNxY/09SNeo2Ddb5dpCICd1Zo0RuO7EKeR/VGIBCKn/lQpnlY3vCNscTAc0JNhIuW5
ZMClIIKjEibz1fEEDM1mZDbn
`protect end_protected
