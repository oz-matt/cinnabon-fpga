// (C) 2001-2016 Intel Corporation. All rights reserved.
// This simulation model contains highly confidential and
// proprietary information of Intel and is being provided
// in accordance with and subject to the protections of the
// applicable Intel Program License Subscription Agreement
// which governs its use and disclosure. Your use of Intel
// Corporation's design tools, logic functions and other
// software and tools, and its AMPP partner logic functions,
// and any output files any of the foregoing (including device
// programming or simulation files), and any associated
// documentation or information are expressly subject to the
// terms and conditions of the Intel Program License Subscription
// Agreement, Intel MegaCore Function License Agreement, or other
// applicable license agreement, including, without limitation,
// that your use is for the sole purpose of simulating designs
// for use exclusively in logic devices manufactured by Intel and sold
// by Intel or its authorized distributors. Please refer to the
// applicable agreement for further details. Intel products and
// services are protected under numerous U.S. and foreign patents,
// maskwork rights, copyrights and other intellectual property laws.
// Intel assumes no responsibility or liability arising out of the
// application or use of this simulation model.
// ACDS 16.1
`pragma protect begin_protected
`pragma protect version = 1
`pragma protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`pragma protect data_method= "aes128-cbc"
`pragma protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`pragma protect key_block encoding= (enctype="base64", line_length= 76, bytes= 256)
b023qSkX0Xle4y9BTjIOoTaNDuPw0OgVl2FZ+nTf4QaVGxdxdj0o6dY74iXg9mAzBsP2LXg8CWMW
dqF6J4LUGnNF+03iIBtho+Y9EREEu8v3hzuCvcuKVH4IqO6eL2ovVzhxVefQJcBOnjPLWWAqO5V3
OQR1y/TpMpDTswBTS7ZnFDs/geKvARX0T0VJBPMbhoCaKVLfhXOAds10tlg2g4qjZNWHXJVilEWN
Bp0HlvZjHGuY2KoAEp4pOm1Qg/sKByLkxi8bq5MxdxEQJ11l7D2uYxNx3S32Q01ym/zpgN2Lo8SR
rDNZ04SC3/H661qCZNWjoWNG/Gvi4b53Ucgpbw==
`pragma protect data_keyowner= "altera", data_keyname= "altera"
`pragma protect data_block encoding= (enctype="base64", line_length= 76, bytes= 11120)
k2L9bEqWwvQ6kZTu90zl3aBuzoWwGKb1Jga2HtdluBgArMzZbv0tNU+8/P7H7TflWgU9qGREAJ4h
dgpYkumXDnTOmAu8jHhCpmS21APESEy8tTOzKH1pYMCuEbkG2gy6xqtcOJ7h2HfpDi4J8dLoqgqh
l7NLjD/gDVs/Rb7cWhCPxtHb2ezkOJXP0rBewJ/a35DLvyWijunwx8COR5mYEgpBwzjYYJkMdvSl
BMF3JG2NUTTJS9FBJ6FFRTOrG/gycPIvUM9hDitLUMLaoylhgNxpu2XO0nWrOb9v56pKNyAatEoC
oFlGM2Ok5TtgmSFd3QySziKNbwjnIr1eN/hmQixtsK1d6zhHoz6tpBBzNbulwEyxaTcj+pa8FiBG
WRYKp51i7QzO+NaV+AIZ5TqsC1qNRoxQWh++VFKqCOhBW8LuddNqBcpSTFEFTY767xEkDokMcf8k
iOludabHs5BGyxev4dAjv3ePibfc1FoCJ+C1xdxKPSQci5V1SOogIRljwB1pUFYz6DgG6t6XuIk1
GuL1vtaT5ynDvse4nmX81eulMsAtIALl6JFkG9QMFoXf5E5/k7MtVBhFgD7/JPOS6hfwddXLK7UJ
diHvc5YQ26RONlGHwuQM0H8VFk80A2XqC7ZLbO6jdGDJND0H4WuoMLeUPEGBouT1izTRHCd0FAqS
ssO7fd3kafUzcd+EiJ9TVbJTMUMcF+I8cwmIZpwVyTdfAfCZ2k7PihbAhyswzrEa9KbrTjtfz7PV
VcUybCDxtz0fRqJeiwyf61r+WPiRnQutd8p9WhpL0QqVAzRm8D2xqamnnxOD4HKekpwVkklHCKOk
PsSEakX4NlQEQp8O2PFGraBjWYOujzWWYyGoeRDw+t/HS2xb5aSczTwLe1V/4zoH6+GTuiWR3X62
Zr7Mo4As/Cov/k+w0JpR1MdZBMaumNwzCUZyPp5ikItnxRvGrXu40XPtzEHuCnMkmN6ll3MVmuZ1
0GWjue7m6AiO41ze/QIXWpJRP3huP5lvmbYLy/seRCkTXpLmR9W+tga6SmK8Sd69WjRfyuz/EkDC
0O4EP5x8KAo3AW9UEOCodP9QpyovhNXzeV7OwX5jjox+PMSVr19elmHwnkS3kAXzIROSyDTpW1OK
3all8/gcGsNojPqQlSSr95pvdFqofihCnrXs78l00YCuBH3S7msxuqPNNY3hN8nmZ6nkojJZvYvc
gp9MUIXeKjuKkjMHCw9MvxaX7hdbURTr29z26XHVupBY/tHZAbjvXz8vYEI4/j6oaSCg3xRJiR3q
Fn/P5u2a/pjDA8NhYq4Qh7yuoXFPwGK3B3qo0ozOSycCWV204zon3rH4buQELk8oWpDBJuz4T/qr
CUa4m0hiosgDX/+w53p+Js1eK3tAVoclmNJQfnSSt/4T4Eba7LEqJ06CCaULPwcj9DexhTJ3oBZr
ihmIdOFuu0g4JU2z/xbIOydWPI2fJvINCVhk8f8HCugjuy8ii6YALQIJDMqapKZjXm0kYn7GEuTv
ENaSRDOEup0UoE4vWFgkKK1g7tw0zFnsGeVDKWtRWUckY96+72Us3NoLW8xITUDhM+aDVUdbb4a4
dyHJJyn+ADtCD0RsVQlDmWGQct1dRHXxU7uYOifG9yTroWVIdPvF9U4ELKehTI5Ff169GBqZyTLK
j9vzQvyvXKmiNRtyv87f+HgG58NQt3l+wKpnTlJsiMs8YGA/kJ3Zdm6fVPVqJ1Mtam8oBeUbhM0E
D4XUjLRbhsxRiSL0NkCoOn7bt9VZqYENZBhTFw26Not9P0q9bOOxTRa0FnW3tWiLX+AsNCt6QjWq
peWXpO4K7DHV0qL9ZxeT8ZfG2Q8MktaQ6SnuaMjgId7Wb32eyFWHXqAWWf7UsvAk/zhUfPtmmng3
bqdLJBzHuKIvqNwcN4HTM8BULGZ9JJjbOalMP646YxLi/Rl8U8mFj5slfn5ZiRfX53q/UVBOy+1p
jXIN7NOSxrqAbqj5rXv3vrV+ibpGmCHKOSnOVvZ+RM+hoVQQVL3gHIgiK5k7UpcQJ3UF6NlYmDoy
5MTb72Tm8oOpyBnq+OydQ91ugC/d1/UDZ6d0+Lk/4qoeLRwGS2hb/NRpmXGPiFATJqrxm+mp6uff
6vnnZqJ00/KOQh1n26xsS7RAqiShkozkYPMQMJLnTJe34A6DMmbtWCrLgG8NrW40InteqCZFKTnh
ggPNGG5u3dIjERG6U0vKhAsIsdoC65prbhSfQuRPeS4JXEs/G5P4hvOwpZvG+/31Psipv8LIjJff
dLFS76bGm0g2Yba11qOSmH2W/kh5pMdEGroSYN4x/on7Pe5vRHS9EVmbrFz7UbxqTz8sp63eEvow
G4sTv7WP97d4iQpFUf25vTUQQNHjIl1a6L1N+wgt+BtpNskqSDPscH1zIaGjx7DlsZrEMxNmy9Tv
lQWt7ar5VdIIsfl/quS1u2YdouZsxq4v/tnbxrmtjivRtQENR+soAnInUGfFE9arBoecViVZkNXx
DuMRSCscMeZvDA90Q5lRyTkjpMfTsIb38o61yeM+kUpGG3Xtfp0Z8YQWsYUYociHzUY9deH0WtHn
O3Nk/Z6klq+BLiVQSktE9IVWDCfAOsWULRv+lF4xXysWrRi8PaWod6I4yTsKnQSy0adO832lXKCD
KLZt0yHHwvzyjsJilFCRhn0tPcbfmfNVlMX/8GDSJXDS9HiS76Mnyyx0kFZnJGE8qcmQUs51FqbW
2XJh3mYcXGiujXLM8wWsWvHmTORhYldrQ5CL+LQJI+A94lxTWmQdUFREtQ3Ql2swY/1MBAkfNlm4
NUVJ+VFYOLriWjyGZxY5241onlUOGeMUCsXvOLg4ZD+s52tu2mEVz93+d+4VEHqbgHBoWGQwDT0r
NEdHOEibxJCOL8a2bXQxUbP2W7MRSFmKGMNStKVvjxG9T9fBm519jl+6yRUGB7IpBXvlybU5Q/uo
kpha2/6JMIHCBmRwQoVsAUDpWEaIzV/fxCtKsKeVagbbkCzUe0vqBmwutzxtELgHhApk2LAxMQI2
mBP4FKYby0gQvjFXiIeSLVDR9U8BbpPrChEy7pbScCvJI3wO1P+JmfvonTzKlBqOGtRv832+n7rt
ZjtgzGeC8E5jRv5ADrI2yC6j8yuMcRpi+s/c1CYjv+uwN+FOqtl0wSFwnCc1ZXIzVHW8E5E6NxiJ
/qoP/f6bx6Ul9SqsEtXNXkSvpZC4xkGObA9D26yWGuuS+542gprdG+JLEG2OZ6bMRRbkD8gH47Ma
O68M1aOXxxORsxaiHOc/fpEDv1pN2SRLDAe7a/YjnC5iXmO2SScX/WU4sv/DnPl+B2YtyP+tMKzp
WBI9P8FXd1JgHWzTSsEWnA1Rxh2bXXpBRLnQeCYwHV49Qo2eI6WyE1wboQ0F0mqyvSXqCU1SinY0
TqDzZZ7XvlK8AllHL0ZW0QJQhy62F/6fPDVEQorGIJ4j8/A1jKOeIYUkZw60QQoVBC/0IEesdUdV
eUMnPdP/RwoTkncWeUR9AOB25RMnDatFXJWWbwlBRrcjZbviHzcJc2OfXnh1lk7dykGbsZCxA3H6
nPPylgWNMwbjm9fdNIPXzb3jv/BN4J1C0XjIQF1W+u2Kemo2xs6sKJUas5z2Bfz4ht1h3G4U2aCE
3XYurDMJgiHtE9y2qgK0Rw0lLBnYrAbNygQcoSVeXLdvHPF4LEhE5Qer+xEj9fTyJUVm+gre6Fsn
s56+Cc3dIwBsQMAUoIrbyBUN+uIFYbvAQJkK4VY3z80yqy4TH0ND22mgYsmfxK31PsXVNNHnEQ3i
dsAaJFbrXMcrUW0bwAZMZbOAqTKz4I+SQd9lygr9kUfx3TczTvjGNmFnkTjQIW8NRnrbZ5f/xhQq
D8wVQSprr0rC1I6VAhFvZXBdLAaEOAjhuQFrB36J+whO9RU9mLXuZhBveI2b/u42u9GenUw0xERa
i6fhUTUnlN7+ZRgFPWtrlCkfjyxPr/ffxWEiU8og2ZPsQDN/tKcN/l9fBCcbEt14sbznU5nVee0J
raQIYq1vEbKNdy3QlYuQN1F05r2ysOlFs47vYKbgoz1mGjdCYK6WZAMomcAUfFeZKBfhT0K4+4z3
bMx4lD+5bgiQQmhW6XdcXQU3Oo7yV6DudVJUHS8KHJxAEEK+q2SraiBUkzCSDGvhFF0uZkUWgJAo
phxz8u0P8/HErU9PaDm+KGQuP2JxI7r4skanoj5XZnZKGlE11uDSG693pltfRFTQt3qXpy4cj9vW
rMVgsBllSvAXpQ9GDGpOeoOu4T/6Qv0zkYbUmyTQ4vIZ8i/h+tBEAHDoNOih1Zj/aYTQvLeuxjui
t1e3wjTraXl2ZQcR0Euw9Y46EV7XqxJqJI0NEUnDrKDx+8CIal4gVOTHKo60muB/v4BIetQo9Kxd
lNDaPBh2hRLqtfic6F8BV5Vwe75XePYnHgCChKzJGF4K8VGnT32H7nB6VV9OiXzYGFWrqFd9GkzG
9DM4Wgu89xFdmikMlw4bZTniCW1+9uFTVHM/jEe2ejtBn4YCLSoX3pbv5TmT65Pp7lYQX/Ti3cnW
3NGN7pOYBQl3JwH4KvHgwEv3nvqcRiou7COzNDYU6P6EGRqyDRkGyPS96sPLRObRY38s8iHisDAO
KXvBzyqDxqCkxuMuZAHgkUhxUEj8AiMVqmqvcINiNqvfjQjyekmFuJF2BJpBmzt4RDY1cQPukADm
8anuwXRJS8ycOtHfIzN7isQiV7NsJYU575abr7WXI+ZwS/39TNTBneqzbzPWcu14kd9byiqh3RPt
J17UKL1/UrcYBCqQ6Os2ItXRBtccKqLGj8pjbs+dHDo+sKmguZ5p5vyN2pAhWCEpHiR2oCWtGMfd
T8btCYQ892DVbA8IiTfVPujWNDe0x0ZDn9cN36RTiRG3y8xo9ta0ss5J8Ju+YSjkbg98mwSWL3L4
Wg1MfbyO0JnZTE2a5kEqgnVR6XXAMpkn14/oIjnehNriVMKqUxNP6o5cUDj3CK60DighEJtHie3I
vrU9H2eZRrza8KgNFzPtzaz62O5+WFOjgpmJN6J0k1BitUMB8g8hoHbad6ylRU4epsyMmY7YAUqR
yCn4QRNTahoZJvdbWW4CLo+0GTSh0VmfW5Ua9bIhIIlXBSgIIhOVdytYljJI6s/8gfxXOcIgj588
RJpOsdATDhn50k11iW98r5bjSE3/TA7vR7o7B1LZ4GNERS4zwfBi508HV3yzPZlASz9myEKiHZPN
ikbLobEIBS07bnPh/yiOlr7ynboAyN/orMslmVWLgKUHB9M6Q9OxZyYude1FwJ5d+qwacryTwvgA
xgvy6o9AoXrEYAlwjvTicEsuutzmoBikvgTMYzhT7I7zZkK9rOby85PkMHWjYD5ztdj38r+sgrvL
fzvbIN7mfeaVry0K68+ZRSOcVRfum8vRMouj3m5mGS8gN6novfujls1xlY/5mVdPCH3IfB1cGAqA
5Y2Puq908E4RDUzX9TuXIPSPyP4HOZvl1DVqXhz7+ufWudtBv3mMXfccIRhL+aYbJGEhmomhm9J1
nG24xdjcBlvxMs4DhZ+wCKv0XC1uBQlJ4QS2671ftXWzGRbD06KL7UpG7rR2JotWmm2KzNJwIaFX
ZqOlOp34Nc2UKziZsz9U386ScAolnJ7wxYvG2wZD8/VKXuURbyVKzhY79cPb6WJK0P6AUxw1lD9L
a+a7oFbiCFmPiFCooghirD57tDOA5x5toEq0v9FhJu/iXZS1NVU7iYFJG7a31EZY1pO8fDlDbkr4
GKIYi1RNyWI8KhkTdNQKdAOsra22cLRwMhE4p3I0mColJ4bGJ5JS7oN0FfoOmTitciyATv0aBxVg
11j+RBZXRJ0TYMndfCtvG4TZhvhLPb44uojwoglZdoN1YaVtNi2KbM77ojxQoR6d9thmaWbsFHvV
fD1oBFmJXmqMQDsrYZ7tIAJEdIR8VNA72DtADJGOEVN//F4ge/Ddtp24w/tbbA4Aiht+rvbdEZ/T
/w6PB7KO9cwKKYakvo6bzmkzw2LkpWcnuFimXAbPMYW/d1RWLP3Rlg46GwKJpxgLeiuOG4CR7/t+
1YfZhTHCmF3X1FvKyb5jKtTDbSPVirrVbtvjHuBeaMqDSAgZYY+dBYqrYfQdkeDIjN7G1bzRMjC9
mZG2oG0DJVAUL5zpBiQTyd8AhOY2AxqqUb0QPTRP8UOVGGXoPqNwO0umhniwiO7ykHIlAeREDzM/
bnXcV8V7fEQ3ERptQWid/JPCdOjs0A3M5CoFNN57AXUX0QEXnKV9A6pLBbloWNMeuPsTqTx85kuS
zqopbdvHdJWPWLqTz3ngb6RfbSRAYApPG8OFV2YKXqeAeCQHi9QQdiZZQ0Lh3Rn9GxenwUyO4KqW
UlubAvJE1u5UcvWAKft6VKVmafaz8xIWtdSJ7u3DThCSqynTd01Z4ajkN7pcEd3a7VGBOQxATxcs
WIkGl4leyq0KZtQwN+AVvDohxmYQ3OoFI2xKT2nLqm9Px4aOwKajN2v/efF+dpElFUxIpPDdAr0b
vFP9NUbwhTh9I4+VFz16mq+PA1CRDnirW4XXJLh5VpWCgCvprqNSuepytZvuGZA7HcrPLtA8khKq
lGjz6ileF9r0dILo9g8I9xRZ5G6qltfTkB1l1Nl5EIl7dxxwZsD0Q1mhYWm4rwp9ckYVSvPJe6eA
rjk1Zjh+Nx2hwKK7JseShFc6qogclQvc7PgxuZ8XYVXscmxwu/rnPrGJKb//suwZP3mPhzkzBluf
K86tTJRIwzQ9RpPCbFp0edrP3x4uSm24Pxg+EF+YZHro369MvVGWlq46YodHr2PoE75eH3ea2OtQ
8amnwpSC0gLML+emlUgMYBDLuKSeILE6XDM8NYeTvJDXFf1wr6Zb34l1jsRdRwx4sRfp1W/+S2QK
Oy4yiRxf9QEowNH/Nfk6XVS1TqA/b9+eGfzRXuwKjAbC7rQ/tXZsdnYBCK/G6t0MDWADsLRCU2N5
4LdMsWvXczQJ8SJfmkJXEi0m+Pwo6txihml97zqT8quGztC5DNey/MRoyr8+QOLMq85C3SdV2t5k
LLBdbJz0zOwBXoMvdnIwbUdKCc+UmdrHLcHxwMLpRrDBIX5VisrlLtRzsHO9W999vuGZcEptp7en
r/rB06OxiFNdwa+9nt4bgYHtv4jhDJ2Kbw99/3k/G29sgbTjmHNMUGP1ThyJHFJFDR1hsYb2EfCB
bBVxtp+sfFKiLNngfGkmAwz3czStJ4gk3itYq5N+86Hg4KsWlUqKW1biPVgm6KBc39AHz3wSDW8U
VYTszcRdR2f2wvrMGDRckt8G7jxvxX9Ze6oq4o4SoAwJ6aJb7GAgHk7zFdpMOGkEt4nBDz+Oe72Y
T/v3i8mxMeEHR/MB3KGR8fBdEVn60vCRGoAOSoEC7C7EQ+uhdBZaYVUrc3qaFf++KonUNKWyX6Bh
4mTJ4YVaoe6/uWYvrmRCQd1FYN4jpyz1VRL+ql4M/ohYj8C71qtXC0UbO4wGNrTE/qi6NOk3ut2+
W2Hn3U4jq8hMN+60hJ+4RH3IL61P/+6lhEiBMBkZFx0QC5a4BOnEBKrRLMeUcvRezUA3O/IYrkAO
ECLFL4HaliMtkRTd2EWwZKXYP1WQjsHUjOVsk48OfexFeQspvtAdr7T+bh9apYnUYE2vM3TV/cIu
3teNuiBWzSNDf9Gd24zhfK552SzrWmQ6KNbRePUATQfbvz+bFNSsL7Uqh0MFWJW1NIim9FAmldkh
Y2xEWo2kVrH+C4m2W8pmVsbD86+p2ZH3LxwwxvWNTfZ11l+Omm5deTmMWjOZRRw0VwaGotC053jj
PyxmjsUhtIprxZamX0om+HYorRvGCOu7DZ0qF8VZKxVl2p5IEgwMdlZRgzgY4u9RD3UDPdEFTm/o
8SdClvB6RVNMO+0MMS0JPzuPFvSNJTPODj2lex1DuSHKxXbxGa8oHpmLmLEAiSkI1VEzdRNyxpcS
tXueOTs8I/dXO4xeZCsVsVHxwKVyTtKonJEEduQWT9kFY2J7tPtzhZ8Ft3ZUx4IjA0o3yz6YYJPb
0yFXQc7SV0WbZrzrgR4mOr9kMozNnpuZsOTbdZqcLDs3Mz5Gg036Y4h49fwpZwCEBANQ23AZXaco
h2nWxJdqTMed91r9j4pl7oqv4j8NYNN6SByLFVrmCfE/BJVygYlYsaFgzb0Qi0761tx7ipRC+Lv4
vVjwssPyJpGC6n3HzVg1nbPO9qDoEQW79XgMaVVKiKJjMR0lfIuZvoazLOnE35rvTCsVIC8rvBqS
mUKvCDYmnXZDPATP9aTxQLvAdhPUUvZXOM1g0JPtJznNFU8RH2tzDemGuR8615R198AhrN1Pnx53
gp1xzevuGk7LzIA55Ov3Ofsg2V16HTId/vWFruhsX9hjx4jFvS7expL+7JgShB0tfTYf/yiAy9MN
Xsh6QtrPecH2zw6UdsHUv2Z+q0ApT0aZHlhvzkNrPLolk3Fp7dB2d/+cQhJ4lEwZRVF0oWdqSToq
nu5tMLlS0WVn90ESkhn0CNvZGhF7vL4wwfelEuduc/ZbLuvz6j6aNiJCBVB1FtzXj/2WRJndc5Cy
Bpm0GHKKOjShGXmJ1Q1QypSV2UPEqomlaypeAM2sO/+gV/wtuZsjcYm3iLJVW+5RGnUEjBgx2FFn
q5wx3S9u3pMVl+eGQhslhPrTuWTXHr94gvW7MLxE4QfRvNjD4uL7Qo949n3vJqsJiMZ0WY3RyfYQ
YVyZSydA6UujEh7TNAsZlEJnFDwhFxjbSUYvizHyNo5WMCQPcBXzDjJZYL149pAwUOZqsZcPWDoC
qtupPFj4FXpxqdTiVeY7Vu/dV39sjIp0ZgvskLzLul6ZGMFWRZW8C1WDpzwSV4+gkze+sriVV09Q
4jGYU3rCFPLjyIDwEefH3NISasJCP9ebuQEe0Fa+JtcO5Sf9ODOUjCdQ45F6MM53dcs1g1nhH/dr
h50U8EqIkzBB5cZFCFdaqwO0rk/a5t2RgS1rn7jI7LmyuXY+7zITPml0zjDxoZMC8PrllsOx6Ze0
xkrE8OYhvLY+p1MyN+4wLcuo1eqvig9ClMNO1/szJwvth+qFaL5+EnPzqv1EcLlbRnAbWxMAGy/b
ddmBZFupChM68RTTwp7HYGRISUGOJPu2VX9OXiAvpmax3Mlg9LHH9aJfkcpj5dXMK1wVMHPTfic1
XQHgrr2GedtLsxTiD2lVob/OtAolFFlGMTSMzWVMIml7m+rN3lfIkZrgPar8lBfXYkaht2rJ7An5
OiJ7GA4stiNpzdIJsS8roRWjbTvpQNt+JGKpOf8d1hJr2o+UwpX8NUXEvjZpJaBxkY5QJT5oPdHy
0hk86EVGXOKj7qE9jnyijIDKI4P7Bo+Hnn2iaYDyH6U54JtwBDpHZFBfKneHObGjm6t2YY+O0yQI
RopSIUcLtEbHpuJFWmYf0E6KA75ce+/RX6uV4WL8WP1O4dO1lYclUplqIkz8nkkjFUZI7KuNmG8m
4DdGCpll5Q64mV6fLpJZtB7aRktm5n9D/wkMEbZt0UC4elgh/Pa0TAjux6vUtVh/wBNzD2jQtzRY
TLgD5QfMsPhIIpYfOKSPEgDsVtEjKbEieiVwGkRb3E0A/lwwhxMnRpkXJChcHqHdElwTVxeAs1vX
ipILWSmuebR7FXiPT3Fpzog3Q0FnMucU68AI5xMmmeI1X7ePeWs3XfDDIOK4v/5J8Ufld73+HFbs
Tp/y9ENBeqQfiSJko9TS8/vG5fKe8JpMxm38xFIXysYfzUfJUh9l+cxXYHvv+aPaAefkb/791CVx
hygYliMUNDMgQ7wt1V2ycnSjlkm2pGd+B0+CktLmRcnDirdTlbSnil6/E7UTosa0rV0jFsjLRLHf
sDK7qoesipzdfbYeT06ke73T8xfD4dth7AI7p39/0dgo22PmoxELq/HRKDJk1fNyL+5aw0BGS8Nw
C5x4KGh7LfkaUGCYrxvfv2rBAvChr90L5BSSftUoPLtjDFOlNkWP43ot+xZWpyPSVU8VQ0X/ALYG
SiOEcv3PjuTPMQZ/gOqqo3EsmP8RkmtYdn1I0PwgqQ68t+62z/gPptF18WAsmb3esOKCI7Znfx16
5GrYsO3LDX45WmUexmOHfzfBRCreWH/M23xgjkYv5eciGjYWQIHJcKIE/o/lyg4lqa/EJwoVFLW6
FGNhvW4pdvZYVDoT+OeEB4opKGsXRHgqyurf3Sc55R3gtbZm30wPv8wgS2WMYuUqCJVjusV6u/FO
mOzOKpP1UVBw1QY4t/riujZTqGMOUV3FpQfnzbavTy7NcaIFCoZhtsQxcEE9KoGZAUs9CKtMVp4z
uRB442bBV7wbm+wR+lfjDfl+8T4L+EYF90RXTbhkf0dYGgfkAeN5NsHjzuzJvzd4xlOT+QxJrSe/
RaEUNxi2DRVyZmeDLKoxtgcCumNUzt1wTTJb1/fEIno8V6+KBX1L99zd8FyGwaxPAuW3EFNh/hXP
Fbyf4Kpazr0EHkrushNEJhC0zg1sy5HwqkelcIe62mX70RJRrh8TWcfxRff+2kfpfBOrRNnGCMf/
RPFBn0J1q9tdGUp5wjPZRrUmwf32HtEBijFR7IXLVqahIgKBg8EuKWUSRTD1A7bfcFkDGU6C/syR
NQ+Tlu2p4Maw28G0xDlSoC0mGU3OnF6m+q1UrWRVdvFUmThkpOkLDdJubwiZSK9Yy/bJNJpnaohc
cNc+AqmyJ5BXH14bPaSrZQf58M3UrccQFRyDXc0LHmqKZGEctizi5xbBFcaedZXtcWIGAumKLNNs
yoZQCgs5Uciok+ZDLaiSznXEGTglC4Z5sFM2f2TLNGy6eF5WdUd+gqHjwdGOx0mEmFYmMTQcMv6F
Rl5MJbYrY2I0PNIhgiNBZYqwIil3PHWiA8EpwHSjoF+co63lePVtVmSQ6Xj1GfUgkGYd2TV+yOhX
ReouVowdDJOKvpVZgpiJRHZW2B/Zug7bX00lD8L0hceUx+Cml84ec7bjH/unKUr6qDrvHLM2o8b/
YTHIQTBJIWA0srFm9s40onqlgF4dxl2joO62nOZiSdnNtYnp/q3QIZWWuW4ivLOsuK7/xNKZRzCL
mOOLrbyw5VD0ISD/U7eW7PXB3k/jC8IxsBD8QgiKrNlJ0Xt9tiVCT+srVZHZGjXkXwUv0vJ72Q66
wlS6jsiLrXsiKpplh1ZJTN2maeDqmvZGkXcmHRB7ZVnZEj4nMFTBdnxYckNlDSz/6yFKRt3qkvRQ
zq9i26vUYCnDgIQ57EGzLHS4usUKpbYLusZM577PlNJHhgGby9SsaJ2TofWNU+FSa1+dpHGdKPbA
zBSts/rPWX2adCH8cP6uCkDgHCCjKJQQV9KK+emC64ma8pbGSD6DuTfeUAcVFi0yjLQh4dD8bySW
x06sT0Etyv3Yxr6GbcjzUT2D6/QBKAXIL37McyLMA/vmVOQilm0mkYYgWnW9WgPzT25TbChXgDu/
d5+QFbVgVynLa+xSAoHnQvyscioTWgykubMJ/vRIh45O4IT1ex3DGf/43kDmbK7nnLm62ybXu0R6
9lQcBd14BqRI83Kor94Q796Ew+aJq5N+z89ZumuMaCBCfQ/iulffJJKR8hwe2L/w9CeWU9zjRWrS
rQnO+fYiexxahkr6CK0KNEbeXXKkdsFGKuyxv1FKK+CnYDBU3JoGNiCvWrx9LGiUlrEmNFPtZpBI
E5HVR0FL7elEJSFiHp7EoUOM6GJRY+Y7DBm9S5Fd4NfKmYSaHhBf9RlFNc0SrskgMMpi37Yq5SOV
OhMLHmDfxkbAkCnRsgRr3jRXGnAcGu6s5RwRMf1NMRWKQReIjE9TXRfef6HSAu4CW5cDUUpx7lH0
R9tOQiJq9G1lqH9bRzog/+Nm4ZfIpPVS+IddKVrsECmO8vFGmT9E4q+wSgB6e/g2moA+StU5dXP1
dg+v8OrOprfGk9Z6eGDc8ifeHIez8u07vVEEarPEPB/v3+DWjIHYsTRaX/gKVjGtpYzq6tEmReWS
rr1MxQxsY7pVp4i5iL3eVLvS/bxKCv0ke5U1nlNvIh/V/n7hkVicyYic+IcrbEhO2jfGHQEcV3t5
Hn4yAyuD/JR84mnNRkhZdMEjyRe/Nhaqsmb+7wyhEieZyaDi7Y5VMnOImxdASi+d1DXNr3KIsjqO
BlS9whsNnvlrDEpQxkdwDQ70B69kWdyHObOCZXnWGhwsKmkqX7V+nARgAf7X2GECy7/S8RMr53mi
MIeZF8w8xPoeamvJ0N54dYoWlbwPOJsOxN+zJ0gsrhtxbmmUg6JT/wBTQASByORHH/4pSmyuec7k
gRH2nK2EUEcmH0YsUrJIiQ5paYssAo0VLlZ+FBLfEvlOva7rZ4ICEsJo/HnB0GQm0YDNLqw59Qnl
etSN470jzzLHrYzqOfwXm6wqs6kHVUm49GWs+VbALqHvyCsuLzyD0QhbsIKIntGGiOD+UqQTiEEa
N9dcPhFkcFNmlyTuVEgkkRdDm0JeUQseq1czhoJwmgI5MfU3w2I9KcH8agHZDJdqLM0etORtIf1j
ykCYDlzwkaqcipFONZA5iF918LBYFrOwud8Rla0uwjAX0JRVJx+TA/PZP/L/yAYMzXJoUsKSMVNG
7DFU+t/WRIMwYZApdM+5MeWotnv1dwy2uv5EeWLAgKyVFnuREnc6MCQW9cR/L+ePG0AeBrgLhEKX
Za9DGY84uLqhz+2l1A9xefPVvwI6w2ZASU0caqUPLXXkaviwMODIsimf7hW0WuTPfKYzVxRGHtd1
j0UP7yzBBNRNueFG3uQVafcpD4Byb5wkGLTQRFFRsTgPZeQsRUHYcvZSbrrDaZdY0u9NXva9RHpV
LzNKIpvPQ5l8ieRxtDWlJzTp1cVee38PId1X8W414NehQkeuJ7pkMXnhq6vKVVhxjyEDD/fCBr26
7ocRtZ+viung7yqTBmYbO1ACCxpDSobqOO79jEa+fIqynnurWISjgatIf6DX+8xucgUB3EtV4nw3
dYk8KVvy1BdfNkGATsxMRpUFSnJqEL2VGi3zxvEUscjynCgQH4yRMTYUfEJinHhZk6fbJf5AljZM
imoqoGPoo89XHGxCgROzkKQEKxCKLkNhftzhWHLto8laxXr+jWLCrGkkLOnoOF8br6hjCke24uph
0UC0sHDL3t9ptmSje0CQdQG2uwLpG4qoyqkcg/vlgLcHDh48FsvLpOc8mPUtRVDquKq6txD1aDIM
FjklnVBwJQtrmDYbywSwIJGCeb3kCLRJ9S1w7MpPOLlDtz8xMbgzeWWWfs94/6GctbzqYXuyalrN
s77KMPOnt+zIdK3Fmon3G37cMYrkykkFn1Ph86hjrAEEek5P0fxOgwQdP4OCyTcHoZ2fd6WDbUGX
U0V5ljdddIMjFbGiJJkmZQs/RcpzeamcCmLEnkGgf1KtwV+EngvV7rx/gH2RC7dJtVXHU3gdTDd5
6Mm6xiU2pwJVF7kv3ibR2swiZLN1S+lZYWqgnZtbWZTFZMrZE1TlvfanwLm3SitO7bggChdKIQLJ
X7mPmxxw+G0vq6hMWWtCYUW3x37XM774ytLSnZzwy1/xjWUvTgdIs2hcbn5ZzOFhU2udoxWkh6gn
8gKufjyJxk1GX946JYgLXFkcuAn8Vbns45VWO1ed5iiaeQ0enyyETBThiczqoLeGpnl95Oyv3juI
OUoCw+oPjDWdCC6qaI/U/B7sdI7hVAYQnARBEynWWuQXV7JLw2VYMrirqf7waIr89gEnymD0R1B+
Tzcz/WS5OKA3iMzE6LTF/1KPXfvIIUyGJl0rO5AfiYP6Od8uR9EjerINr9YAVv/a02gC2B7fmytJ
tfB8R/E8LCXJqEkMEJFTiHt+/RzAGlh5MZOJJtwL0PDVVB2MOccueWMs3/NXDKz3unX8pOfls2CV
TQxpq51fDGaTOmZMYXasBQ8FGVqg4TFJxKIdQYIwO3s+1PBeH7fUejfStgy3uEV9k8aryINEGUpm
usvQnI5rEjfyJkobXm9wz0UuUsjrLNA/5g478+iFJ8Q9wop9Wf2HAGr6SuMKWnz/RoCbGA7BR2lB
lzQ21Is86aRsNmrbyi+G2uRJobxukY5WUoRw/iBFRu+t/E7TIXJFzSA43DXLMOMbhNcHfqD2L2cZ
bfOGIlNYXtf0VOB2DOcLFOYHthYhr9vujR7wz0FdJrSRZs6+eP8kcXuqn+azx/0Od85FYiRj3wjc
0HyJETvEjsHLtaAKhPUEIlBXir4a9xJNMgib9CRY0nZ0+Qya6qahJ9KS93HaEpri3uevCkCfNX39
uCfs7JZvAGZxHJIsMVSgMcQJuu/bdyyd5PgmzYAVRAXfesLYi9p6yGt+gnWZjtoQmH5EhvagOiYn
KQ6C3+N5Qv3TQPSBR6Cy711YRU/xQgv/YwdB8zXIE4BikVrp+Ax2VKMLJ0+HiuZGmXLmkgkp/KkH
qvX/sRgHJgzmqK/EHGattnzCAK4wJ5Yh6wwdDdIXu2J+Cf4ZL3tbuJvAYA9cRU29UVVRImlsvL18
H1i5PgPYsqyy0LfYYmC98OJeQNcT2p3cJRZ/ciWXbPTXzkq88b32H7LSREQ6jcZYbd4bcppB0wII
X3UvdF5qY9U9rB18te8JpolE5m+LEEEaHWFm4MMxKo1+SNofXYYQL9Sm6zBabRBkwCV5mLn3l80L
AmX7RStUvgtYAM149NhlXu8ace3bE8on9Mj8DMYBTJ2d5TiYqXDzKz98NQKSojcSkpDfZS7QP4i2
GX4EFtfQyGXIjI3Mn1mU3Ms9lzli8GpISO+kgLXeUgYAxNlS6VtWLJnSDumZmJidDJY48ZEaaDGI
ETP0IAM=
`pragma protect end_protected
