-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VnLcMTjfA/7QclWOXC9E49ayvFHxgskh0naCG8xgcDi69ZYxryZ6F8NE59aO/vJL3RgR0N+i5hUC
CZVX1yLEx66mFI5arqaYI89SRxUWS14kDdhXfxMuaU/+fHS9BlOhF3VXCyDka8/OmjsBTd/ur3Fl
qb9iFD7tNa0fXgIW05tMQ0/nqHchaoFkPemxMObEXy6z/+sYEc64aWzSIVasJEgnxLW2RR/NSnhG
qw19B9REs3UI6kb0pb4uuAaJ9E/NTBlwumCRCH5oj4pl+T7aVJPsiz6Sf9teL3IYXA7fQGOXK6Td
/ssuqoQFIOBplRzkqUQWeDrrN8AXlOnH/Sd5CQ==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 10544)
`protect data_block
XtKcWj51CyTuAysavDvpz/1Qh8eg16syBJXmlxtbhEgz60oTxneXq245rImjeA5MFu69fWf1Rw+T
4cygMqaSuvav6j+P89vrYn8ht+nI/MFAefnZlP0ejX3JiogAZrk9QXJPH7nlVUODBSQVQcC50J8N
1s/LcS/61z2aTT/FjBstK/osYNQgEVbeonQltIXFN5aEn1ZqR0bXnXJOCn69j8q01VDXlpe1jALP
L0/ZeewQ0YO6QNqYHo794VdKfLy6owFBq8W103w+BpkRUn1m+9rlmFjiynNAgkyR8Kwzid1RVdAt
usTHTRS1nMkxlbDTEInb7wf8vTBQR3ehV1YNW/NRYZfhXF2HQC6GDeyreN/ixNdn+o3hVy2Uc1vK
3sgNwNQjzcn+tV/U1Ot1BwjdgTeRMU2AGA+SF9YTu9RF87KQncXzGiEJjJQhaiPtmSk6ZukTQ5QF
vMuoK0JFsLKZ4pOvF3OYzTJsRd4Z/cePHzgiH/RbCdsNjRiWGWVEX/H14byF+eZ6B9iMadcSsEAi
9dfZByVlWL/RzlCzyMOCdRUN7JNCZH4u3VD2z/XbY5Mz00anouEHDd+u/rJW0pSWgOPZDoG5cQzq
/cIzwKqHwbARrf3GbENAU9WDT2GomGdBKqMjiPHclVzfa/t9x5XIgJ/MPlAWooTcxAVLHywqHyus
dc/kFXKcZj5yhT9v0nlYK8YM7tqmPrpgYU2QMujxZoDGRQI+9u/kbA8K/13HAAKqWYcA4UI863Vr
T9Bg30qmlBE2g1g/lhZdyYyWPAZkyr153xVZYEcYWy9pu15qZTHlGMCUAelTXrv0Me/2kkS7gyp1
7xpyKZETOQZwiH5h9J9Xo3p1JPzDuOa0i2C/wRgbdpdJgDny4IIj7TIX6hEXMTkop1F2+QrSyB81
STtnBJiWHnWp03ziZFljCAJckY+VnhWhCbvYJufcFpc3iEIx7tTAsC/biHCahPXrjAyUnTVyK27Y
9KvsdmiTKrjf61mEw6sbJdRcHXwv1qjHmqeOAEQuBST+JNTZmaBML6PkmoOU+DiWWKFsue24QdvU
AaXLSowfzAksydbPTurjz1J6m2tnsJg6OnUa5+awBTe5v9j2AIpm+/z1fVvCCyDBYsvWK/SLSvV7
hPwW/mAZmbHiOzNAsRCxNG5mkYRrdbaSYDLx9LnsuNIsxEWWKIDCL03Ocn/k1aJYzYxm7coMUDR/
kLp5zu/e9CKTXIXdT1X9vGWAE4XR7Y+pPyEKPTEc1rMwexkvVrVDJz0QEnABN6hjyQFkTL+aI7Wy
bBFqceO1C5bbGIoS6a7EpPhixWzewn2yKGaUzY1kQHKJtWSTV8EzvE6sPorlbSuBN1UYXGdQ5P6l
iB/rU79Qx7Hr8y1yKCvzVvbFbzutMF5uE1Sqa2ST0dXKYsJhL9z/r8GhhZpPDhoqN8rqLWhwo+IF
8aXNvr/KiOhI/Kj7SStHCYy4wEEwKMOg2Tdbr6cdukoRecdTgfMbqIKPZ2PUf/JyxYNKhqqF8CJe
8aFK245w3MtWMrcPcE2Vw9IRRSEzb6RiUiPMSXo8UjtKmyjiPMCL9jb86DX8pTuGk7BprC9UqH/u
Mplt2Vv4bq8PVhpArdLxVxb7oIV9XKOBsqxQ+oNb+nmayovyG+/Jbx5amU7HoPs6z2HnNIzoNVmp
cqoDsUBrHcii3EUUG1+OjOFbXuidrfNHYF2ExFMOnr4n3EwBk6TQ5QqSryfis8CZIzbBbrNLI3ij
XHQZjVOAZTRpheFtToPuajbamIZXImfaK5Yyzzhqt7OawhOJzRZ9+TApPS89vh+RV/1ka7t2yF9h
lU90YXZP91ay/5oV9U4jvNGxuxy+WiaR11fSgY/McII+0a+DWmzMidK0qgI2F9jLiBE2cojZqkl6
31C9GsDC3rOJp6zhgmfoB7WiSb8Lx6tRRuXv/swpZn39Kf9n9w3BdOTG96TXwff6qNvcmQWDMtqO
82qRf0MyYeBMPbDbrNx4LEIiFsC1ATKoQiSfO2hCPSz3kYLRFz6BdLy6OigG9zObVrMnjEY0HyzP
07+0/iNEa+l/A8SJPoDj4YaX33pvuaemnLpguwylzydj1Lc+wvUsl74eH6rnrpyNM9w8Nv8OOPg1
knUVh+YF8Z6m/RYh7XGOMGhpPxjryClybYLYV2k+BIdzmOclTxZaqHcT5On19lrtfTOF1aeiTka9
nlB1CzStJ/cbJgCNbpGKIzSzEms8cvWZR/xjTBp/v/GpCus7oDe/EOrQ69YbMkH+HcLnq+1Sy2/8
6qd0EhFjphiJgP7A4Lvg/+BQ5vTpeqpCtQ140cYn6Dd30YMsgBVVspjxTnmKYKm35pr6sCuvjw+k
g+aGim1oO5MdKerdB+NvJXw156cUoJXOsC0UFuQDeozlJWLyKy/CGmOeW8wRP0aVl8iIbNp1YpzY
UyJZL/2RidD2lrxDoMNPYEIGqddgbHwQz0VTP9ijy3QmG34MNrMhkGbW1grt1N20DCcFZljWRUGA
DBRi3NqphS6OoyGl5uSPvin4hWSjF+J004xq9LjXZ0ZzlZIniik3/Aevw4TRPy17G2i2FhYAD0oT
UJKj2KHSnfqjD81ocFAcVrDLS0RY4ZjX+czuHapwl7pUqUNBCvEZVwTPFH3tnFACvz8JI4Zv6HWy
36x73tPyCBDBQAAFKrG35vaGZ9tVBypASJT4LS4re66D9KBXwMjNYD+fXQDt13E5Q4xdBUv4K1u1
qP2gTyHub2BfEnkENxBlSdm6bHq/cVklky9e6rmdi8M6QkN7COQYTIVk91y8N5g47NxU59uhPTiF
MG2nwxJXHP44Rq0wJXeAGeKBDOeMzAb7RyGD8VDnAIWPH88wHXdiMNkHOgsr1dusDSeVQld7Jg6o
n/H9Tzo5K4p3f/howhw5Uq+IET+r8fb66NsvBsu/LUFP2kpRIUwPa7lEKbdkqKtvCCI4M68urYw4
RowKTpoIP9mFAuVl9rzfRZO2MvcKMEPIqVAXiI9QaDBBb4bHQ2vDkuCON7JnQ9XSXSjvS8AFOmfY
UtO5xRPxmy0nYNGzraUQ5Fv+7QDrJ3k9BDiT5+NTIwrcZ0yg06uWxlQBrBlQi7GOt1CjUc4UW9oL
irRkONfGKT3OztDWT8E6PtoPiEkcHhZdNumlgUotpwOPjXnhq2EKsgydgbq1Snok/KTLQguBt5vs
1gL43OmdvtSZ0A/+GpLRp6MAecmPLM4jaxMt2BS25yyycaK3OzYfX/WM/jIXXghO8QjZ/Pp4thR+
JcA6oVd/5r4YEtuvLhWh3gAY7JO21rWtC9JST0d4gvc1IYEpmvFd0tTscJSI2EJJeMjMfWXDmXLx
gDn7X0CRzY0bvKY2NZ+QPqkh9VxHHFRAlzz+jwGCFrNBmFm+AIa1zAhDoLcAbTc1dJtT0JOmGg4K
3HTO0YZLn5GgzE79rThqEMncBXRdFg2cp57z76OxvfEe+eKAzvcvEMzQUkCAPcBb2G+rJrFX5nSx
sg4e9pzBNH0LDu1nBPXfvBCTh4twxCPa8kfOBKrxDqyWPQveYha9IJTM7c4vjoQHIPixV/3pKp5D
LV0wNVt9/FrvZK47tfA9gzERd6KTlgxg5Mlttz1Bhboqu6MxCQrtHnbkDGmxFnmWXP2xni1srJ35
x6fTdSG6NGt1yhKTBY0FbfcgTj6t7OLUPsSGhM3VzTkKYfL9/vSLdcl9LvpmCrkJZklDR/lIAVIt
YrjuEjRTM8Wkr1q3iKxqtV1XnJ/Cxcw1pVrG4pSNF+85nEnmDPeSRi7nwNoQyCgW4tkDAaVj2vz1
TCYHdmNlkTR9P8wHg3sh18/GPzbSYBrgRfd0zMG+7DFcvojkQ+1C2sE8HTuiXfzf8YSRxYniaL2S
J2Vnjevkbqv9OtCswEkxufzA55dAWhd9sDyQ8hhn0Jl81s8fp8tc3CdqlGuRSo0LoquJrWFtcQg/
FhBi0Hf3S/b/kAEMJrW8W3Cz89n85RH+B5UspFWGA+ucby8lJQN+kDnYowyASAk99VVd0NndH4Rk
F3NdUuuEhFSjGRptH8DeXL0WJ0TVcHE0qS42fqHr+Zf3CLOmgNnbu/0No2HJqqWcAwvJGEnQVMoo
i058usbpukH8u/dA3ZCs0SvFKUpAB4fUC6Ya1W4JUWTaSOJeb634kdSrmHPn0PH/+lrb7lbiJA6R
LDnaOB/NMg43tT7FwvbGvc9sEkSYFo+rieYhNITJD0WQCkvFMEVuvv/kGUh0VDDOCCITVqB6s3G8
X7mki1WPxXBuveg8068O6tqb3132egNmwRJgHwr76GHa11qUhaK8XACKTSoqXdsdOsrXKhn/xD8h
aDeJuO2xZ95+a6LApOA+A+YgzNmppEUawJM2AOEuHRUcvI7jh0hat8ZwF87XGAp6jaFkxTfSBFcB
MJvvXSOyHgzuVyyhYnuXtvanmVHVxB44y6+XCTCNAnGSkhPeeO05X5Sfd1M6ejFHlhKbwLoNRZJP
Zj9WK+UZhH822luHELBjnaTSAVVKDknsOWAgKKU0ZKOop7bWt40VDaMTj8NwvZuGqn2dwj7w3aED
kWUgznmKUPuuw/3ylukeA+0JtOHY65tzBrQjEThxDgbwKO9YnCyj/ATxxi/b5AMinm/pts8iPSr0
GHxQuM3xMQr/Xrt8uj5ndRJLh9ufUyHFI9D9Ea1NL40T032SqvlR/YcfCh3ZldwXqawkh9LEZL3W
4YFNRg4CZTwtDTfG3DZuEtKy4Rvd/kYvLnYZR0iKiK/FxP/LDD/+YVqL9120eivBN+sQ4XggR6C8
64FbN/B8Us8QoAHdPw7UBKYWdblu7dT3TZllNdRHG+Q+U6sL+VlsOtxQ0a2gCYRy/q7GoNMaLGeF
KsM1jZDz7wvO76HK6S4BR7ZUfDHT+mSasMpshJf3c+YmvNg8aAFG2tmrx/BPdtTXwTE1mgLoHCOU
vdrLiO/yBIbYlzxuuqeFZ6t3cKgLfIf/KeQejydG4e3PbSXKhP6uiclvHu6rlCfh3Zf33WbokaRL
Ol+lG2FBuKubGCwQOgskHGg18HpBRCSAhnTMw/sYhDPhLmup59gGSJwRN70DzGj+PeKkL7AerzVk
w8JV1GEeBCwngP879saK1r5ewcffXZWzQ4/FyVWLImTczIy5ZL+OjE1ejg8utmhL0/IEgbPLaEu8
x+nd39ZwYGMSEw/1yvlXN8HpD6SnQXoG2xfB1mfvVTL07HhlR/hmMXnPtHAdVht0jiEjFEBQhvSd
762oos0uIrGNliEamYgIfwfKg1SGEOb0bm/bs6JlOejB0FFFy/J76k0wNjCwJIeRaKG3fafSnJQp
n96xPn+4Da9xmhNffC3V0cS0G1YWj+jHqFHIsMQiB28LHukItcs4IKU+xo+xbpYLgxvvl/3f/H67
Z21rAhH55sM44hkeA4ysbKJjsoRvE/CoY6a89HFgpvsGvNSbHSWSmdz33lsXhlPsfFQxbZ5SPzLc
JX0IpjPu16OV4dGOCi+DrP2l76SReMRntkmEQGzawVDmQzPr/0DLEQK7hNz29WjHPfe/3nwIGmIY
Y9lhmuMWrBSLNa5ZHPXJqhEEfgwWZYP7e+mYkYB591h7EAC6Nkm9855Lgd2g+s4G6/7S+mYk71cM
IYYEVNe4hUxhW855vjkJmHr82gjDA2XzgbOWvOGXbXpn9+Ww03Qz/LASXuhpogcAiUudV71TUjUK
j9C81xqIyzFl5PwUNnFJBfH8btvsFh0NlZ8s1N0wGsM6tO+VMSgTYaZzBPnuNuT2mzedA8a0HPzm
mhTZcXn3vksoafp3XC86ev3r8OfYD2dHlOfHTAR2vG9/aTet5v2Ms58HJt1PTy5tEOVVyG+dAmcZ
mPcCclld6RzMgu/WBrCBq/0yPJZKqoyIgL+W3K2ENTRpep806COyoIf7kqA1o1kr/kgO18vFLaib
RuVRZltNrfc2tqb3xO327H+bM0xcGERSzgOq0xXoOnZuLOwh3aigq7+u7Nn2M9kzdkQmYkscPsAh
SKZx2uvDScCo8F7r5ket0EshWADw7Dzod9J6KvC4U452KeToPS0HNE4tMbrxGi3T6dTkAEcXDhW/
I4wbVTNEYiaLjALkDDUG6+y2s24Vdq3Lprd6c0SypSiCPEn8Rc09PooFmOKORuXofkyHcKHC2XaN
dx3fGMcp3s7f+glVSqPpeIwrqFx9TtXIY5NfLJvMbVrBV0Q/F9gp1UbGzpXAvkBHDftQudqkocxD
S82RWcdxD65bQfsrLQ6eDLYXE9LOMWRMA6NDip3wL8vqAmJnTvU/U3Up/DgTXMKnrhbx0xAkDxeG
psM7x6K534TBMxZWkaG/Rei4EVbL4xm6JMEmW2aJT93WCFBbhwLxQTajxwxEZlinyArBrXKomRAd
XsJKLLqSqQ+OT/+FUYAcNV6nNuCvVAbAcr+yixzPrFrqCBSMoZZAlV75KCqw4h7XAXsxtKpxeSF5
uyjj2BLqaaZK1bH7haHmhkYTFJKQhmt0OROp65LeN6PdeeGTmOg93RSiACEORuJD+PhkOHBIUY36
usvn0T7K7K27umv+H8qcaf7E65MvN+Gb6qZ9qpNQgsL93LOH3A5NExj+dzp6lsSGj6Vgq6unjOeG
yM7MGjWDPYGuFTbzkun2ge68c4aLmLCSZ33/NBRqQawjAM+/Ph7KWJk58ZsN88dZ4OCeaB27bgL3
atIs3h/QQjinmgPRHZ+OvbVz+VPKHLvWD+J6MDMrFknqT4D5+NiAQYotfUuKKMi2SGXQwew8xVii
FaRhglGr8CWNckrQETKm6FnW1raSuSybqIqaAurG/+Ji6vz5syzfuKXyF1Kc58dltF4jUKmvD+/c
CDIQvTN/MQm/4jEBNo4qOoXt+yTRV7Yiu/T2EGeZE4hPeO193uj3Sf18eB40I7zXkBPSc2mrwgcM
Opq07+xz6MShxtxe7Me5clNqSggfHYM5puJQaAJIBUzdUouVhDqRgBu3tSwA9U/eRATLXJveFdrk
ZvnQYGW2+cqqN4adI/Hjtz9TQEyF/lSLNGiZs2HpZSLCPoWPHLYmjQk9ffjeFhIG4lpungfA/a5I
SdWqrJ9LM6M7juYJOBfLbNSN2W5wA2dMutiwurboPm5bm60WxY8aDUvkEzVTQ0FNJP4r/GG2S64G
3zJhpezMvDDKaZMa4lFccFH446PlWmUWSn557SauJ0daSebfazydunBnSjDBN/KDNtpPR5Fi/aNI
1SVFP0Yofe0delrxr75Qx24Nhl0UDLEgG90Tz5tAe7DJd+B645Ei+Pbocmrrp7ZE8lyzOuvaIOM+
qzWgIUyvqdpdNWW0UWhNvAH78YdbHqg+DRJ7YP3Plm6yz64MjoZp9CSp5e0jY+K1CIuXBwGhK1Sr
tslJQTrURONrNN1EXJxzDDpGB8fktzCm2/o4oKwXJFwq9qTCdmkDRkci/iN31WaPRC86cvpu4oeH
vnIfsQPa+OONX8fRkLaEXKxNDM3kIy1uJhR44O9WuOKLpdHYaO8IkNBYk5gRk7JK91nf98v/Zv4v
bUV+fQBN12ZH7m+BfKB8oF0LV5XqCEGgQBwFJv6IxSpUWMEs00cqgs29dVw1ijB89nciguboR2jn
n5J/itXd3u0a78eWNbtxZ24uRRTA9ud+yiswNCrtPth+wf/gR6DZw5/nfLjfVJFDQxnSQ29Jd2Vg
8wwiKno+fJkmWD/emjvFlXqqld5jN9Ze15uMJ4zZ8a/I4oe7knuCT00WrQIFnsJfPj3F16fEa+h0
2edcmnSOiRywmo5rXn8mZfyyI4Fw4Ww0VLhTLcmrIwWpV3KydH7tcRcwapRKtd4aySMuMXdiRgyq
4r3A4di1MHk1G4a4fHvhs6tSO/uwmsTycSwngMicJIIRkAE5n/3HDpDqaPbLqnc6S9jhtk2n8RR1
KHkDR2sQloKvfUYeFINptmyqQ/nZnUU5to3T+p8VPUq7Zy9AzqX8ZrYeOwceKiM2abXv1wY7mRQI
2esT8smoRh1ZDeGMFPC+fonZbJhC/Px6aOC0kdDZYQS3XPYvcFnNxTsMsIgjPgv2SyOonfd+O3Yj
StuRipHbETxrY++cdbCp7HOMjAjyP4JMNl5j69QwkTNRMiggTHcXaN2dOH5ocxd7ecxvAXjbvbj/
mE8fesoWSxzyxY7+h3Mv6oAld6EFlAa2A/I2IUvv2GZ/FeRzxDvQLxLVbXmpkxxR3DtIa03pieEi
rkQZZWQWrbpHPy9dIk5Lkham3vnJt6GlSGdEO632x3Nv1npsxpUtLN/f5r3avJmA6TAqAfcnxE0E
yntUNfzuaD20t6U4GdiMRzx9h5iq8gKUrsLc7VI4MSqh2Me8HwvZ/OWBou8uUbArHmoVm89tmb73
WFkm5bXWnHhHLHJO+d0IXSodU7rsgUmghsZt+8NNXeU8wcdAON2mzjYauf0W+MaBPn56Zfo5ugnO
jZH3cMU0/Q2iKmGwfUnf9RBCbfI7/8n+9hOUZoRWjav9im+6WCcZBQ8nBn1oZXC6RltNxUrCkJbr
9CP/haC/C+Tqub0bveHKYqaH1dk/ZBbeFoyRAVjyxoP7xowNC6cQSBZAhLvfwMc7f24PdzCt5if5
AggWnHQb74EKeSJvHSo3y+J9ZcxRHAV2K5nYKDaRCtudpRyX97OwtVVFw5qdcEt4hQwPiSLLOTQ+
C4nB5LJU4YuBD4TR+8M08p2IAkOx+H0+2yjmglJGzvzLWL3Mt7XxhISiQzKtvz9i3wn3r3dshEEB
p10u4w8whqguQYxH+rkEcqKls1lv64nWXUXtzRTUSBaCHEUyVNNdt7uWeMbFJuge5RfjeV8LpDu1
E748Cc6VjlupnsN5zYzD1YHUb5qehP2P1Z7RXGS2kfjJ6wGwTpvX05dVC0G9sNIq+iDbEk9OTQJ4
oSaKWaSzcMWL1Bkp2Y2w9MOCOBaoIRBz6KU1o3AY5h+wP6gK/oSxmfqdeTfO3FFsLLKLp9X+pe0c
j0bAYDsiW09aJzD0tnEylP/xTNY0NUgGQdt1MaZTs+Kc5F2IvHDl+cQ39oIb4OepGYmMzqmljfts
lLViCo62kQgHWBJ2Av0w/RBDWa/8WLKh/NCN9zkU+REVNpyvHj1r7+D/EXXXbENao5YUkCY0ouZO
7hCSO9wX8La8K94BiONYsmnk7J0FoFJqVSdHep1+SnTue3NrJHxvLiihrQJmAnQyzxNOZsd2KWJZ
tWcYNWGaPUgKI88aUFJ2FFNVVcVAob+mCXUOTtLJMvabqDFyp7wmPKouConmckPcGXEi/Mlcictn
kj7Hib824epbzuof60K7j9r0GaiI3oUL4X0BPMC1SQfNcpqJqPgbDRDe/N63ZjfKvac+J4FT/WzJ
4o7u9ixoPsHaWFRdpTvbiRkS4I6bmR7zcZCEmL+zs8Bf19L0x3Jr5XJ6PqCmI1G3OVp64n9hTkYr
0cMFKi/AvzcXb+11GjuWwWpesyrJXPxzjFaB+YhnA2ESLunl/OzEF8OWh5CbZg+9E6wVcpYpwnoK
dIGXB/xxzo35/lRm2Di6rvJoBXZbFkwYDsL5mOUXk4v1riCVRCAbDHER5LuJYcDpNGtNfP8OT397
2VsuXO7BYsI7nzDM/egvA04cqJwhv5QzHJ5RP0B2Wy3DEkrxYwwAY0lUryJ5OqAku9NRqnHi59mY
qCFV6PQnyW3WynVOTVw9Pu9TGiQ+g+mGM4yh1OBB/VceZ71ePvey3a5CpnagJW6cUtoDu7c4L6up
mKqIIGPhFYIxJ8gko4rrE17O0J8IemeCDOp678fZcQM0I47hIqlRr3r4Abe988V0ZL3039TWLiEw
RAm/WCrWYQK/ZDfl5KyCfLgv5iUiAmxBGYeGbgUeqPmsUjIkx4I5nJYEG+AQuBnX8nvXoNUzhT9G
OrpD8GP2mbc5Xu9Mm/44rPy4ic+ySbSPE0So7DNdF4gc/pQzPy1gxesHdu7EDrV945fIkRj0p7LT
QNLefDMUOPpmaNd8lLuS4m7zkiF89GpHcq5Jk9E657Y8t6nq0KcNuaO0HapQghPafyj1NA+lcFWv
H45VZUi79rb1ZU9+9LnDwESaAPYnC+rGglkhVySxegpWoOl1F83ZRBaV5gu/fqU1WXQ0C/AxEL/h
wHUz+A+2/FyWZGVPrvucNdR4h+sI4uvPvXfT261R+psgsed8ht3cCBX0dqlIqp9RqcwsLO3CeGH3
SZtyyONdjBnknGRiYyo4pTE7qkg9YDM/Uozy6bTseJijVkIpJUyw28/wDOJjcBqwueVDSMrwgedD
6WjpcA/ywqXwxJRfttbooeCPMdTbBi+5RyTfNyZ2HP5ZwdP5EK2wQFLul5DqbJVgK2Mqj9L6YeTy
jxkHziR+Z6V8SL62nvahNm/MGVMT4NZ5CE8l2ZJRtQcHcUn8BBSNJ8G4n5Ob/kBADeDYhHlNqDPJ
JZWEQUVvCRayLNdcVevcFCX4IhXqjABLYd4YvQM3TZ+ntWGE1PDTecVG6q4i0xhCEBs2Cw5p20NN
lmIiFCsZ2r2P7eaKrBEge4laNZd40gFm3seHeRNJwH7do2T+8U3HWk9JwBKW7LRkudrfUVYrIc0t
SgA0nWnEAh7SFK6IruTM3FE4o8pWLUQ3qko4Byk9MbvFaBgPjCn9otoDL0kRwexLrdB+xP7lJsD8
1J9VWcVvaQmTUAuAzOXPwNEq61pbTrWRN+E+ROQ97yQyHcZxpl2yAwk/FGtOGdCu3p6wxe/g8HH8
lvu+OFmZjB6sxtzrHj2U8BtM7xPpopXOJ8oG3J26CIUfDlMaIabUHmGiW7lIfSkso56Bpru3ZExe
FHHjZcnkb6JTMlW3zARmbTagN0eMHKsH9OYdWU8Ewbb3wv3pcAraEsN5eb4nCAuMMA55rRIMaQ5J
rTngEwGbxuK/vfIDh8HYUdE4hvQHQcsSKJnfJpMN8zl7/igG5w8QenhV9K9ArgY1iMPAxrtsGAhd
EHjyvJJUngRos8qg2ApwoFGZh8gYMCkUq28iml/CydO+QbdFKkS9LpaxL9ffi1s5H0z/FE6sDSgP
v+iqE52pzCvFyEPMPM+3PfyBSLJj+a11MAbTjD7vyXWcqgNhL6KW3tE9yhUWgSyVXHHkzFxcqYcX
qBvvuDyT8I0Q0/5+eJrEbIFraziBbyZ1mpLbgBP+3Y5qSI8YdPh8YGlBxGOhSw+1gC0VeIyJsGn5
6vpqP09EjhFVzobJvR0uJpcdhieMKssl6wGkaeoJ+kmJ3C8XfX6RxAGTXDKA4TYm8s+ksqZwJNo/
kU+uLMbhD4HRiYhOMODuA4LQNDvxhtjxzMXky0ub80gDFr2jf/VXX3lM5Ip13QtEu4gx6888ht1F
777Ep2ASJ0vPGTtgeBQKZMlYCTKfkJuAZs8dIFN5iA2l0ODwf62pMbDWWfzllz2DR1mxAFfAkZID
HKG2NLEbGeRW65DylJ9swPeefi7v0FPfmBEv1Ql6ocUh5jY8Py/02xslr3YH+2d1ngSj0k/Oxi0O
V/DuWqSBEc5Nxq+5jEYQr1vMO4E377Iem1KCSr8XYblSgTEiN5sB6XJ75tYNUoT+ocmtX/jppfnA
1gHfPzQUjhTuDIiDjTYHFYjkirVHtObotV1UDIyG5BD83/oVkYdcTXP5cOwszy8MCsaoHiuszAWw
PQQIL8fNnyPUrWn+oCgWIW2Fc5FmuEVJ9qzZjQTgAlNA42BVbCQtlyAtyopTdhIX+YHquOK/yDNi
fvcVS6hKg3qd7bVe448loRK4Vua57FBhD36CmTp4IYpuEwMsR2enwudOhMvSwtWBNXQMOFzN/hRe
Skmxs2ocP5lKff3FVNBmn9ja1zTTxZketsvoFHj8EdivzBNyE244sIYZgYC2UhyK9TGfggBbTHoR
P7QIKSbLnURfoMIkYshZmp++sQnKO9oCzyPdcIPjGC/C3suh4xxO4a8C7LCYngU4sVE/AQn6AAlK
5clzpNnKG+8GXWGzj6yrh3sq7vH7H4bh99sAHZ82nmGOoeLGgWSpFeqjZpfDiVGOkKCAI0hTJHU5
k8qBM9BE42ToIC7GigMAjR/lX7Bcb2hMHp479Y2IT2UpjKe0c5VGTOZXgagYMb8xOm6ilq9ZXnSz
6tbYxQVzFdHwlpe1xBxeGB4HuSS3HI3yS+WjPHxim493qMqPzoB97yKRXLCNeuRrbN8pQaj7FBu/
qZgmcNPKEhyAzgejCByzdYvCQfr1/Ln1XgbIyIvlNcvH4BgntYsqWcx/sCDzBKJ8AtLlBcbzE81R
JcPxg8Fe4rGdEikxUhYrl+Lu9FeodF987PuR9y9koawsnJj7GgO6B4ImTVz6aX6QJ90ip58hFpiB
KaGnWMjJcQN/eRKXdq7fEl7ynZUQ6v05GOEpvVoTlwAuhhJcYQUdV1hER2tODva/A1iu0Zyom3L7
FLrrdU2c01vGEWQpTWC/qU2EqKF2uYz6y1EuE1ZrLh6PzFPU0VafFIS8IUVF6A3eWcr0pJLS0GK8
KThGj3egGs75GhXBqVJ98JTlqB18o1ujVYhaOzZ56hfT3JikrWzX93yetMx8lwFwREJNvFYGSYdb
yKe5YRbzOwKO7KzhpUC91xhtkY+iOthlCQsPZIMcur8/q2FPbiD8PV+WhbeCjEEzX77yhQ/bbjqX
7f3vy/Y+vU9XMiEAe/0Okm9JgxLdbrLXhPJtrXD8W1c8LvIZRu4p4bEhWaR5lACAnRirTVaGnW3M
41dmxh1xl8+Lk1e//DOIgsZybavxEUU4X3gONJhLmLcj+IyN9MK82nO41Lt5od0zvpbKER3C4Kme
iVjxPBZHxpmAwyqAuTMhiiUW6RmxPpG5ksGXTvNV1Uk4dTdNpf/nGhkrjBbaMMxTxD27bxOIO8kR
cm+/v3JUp1cmTd0mJktMTE0FI0i2e7AQiv6146zJqm+CdDQveBeG5grJTJFGzZKT/bEFB0oQBwkv
hbc+TPccqfgfjGsaBMJsw9VtclVQmafi0vQx+9fcIC1yinc5EG9azseE9HedH0LJ7F1E5CT6/nsG
WkxhNhgQfi2jZ79jaLACGkRtJImziCzXMs1hXz78HYEEgy/SQA++6ha90aq3Eyjr+Wm2vQhQeBhM
bi2kLCmmk+n9I3SJSj+FIl6dI8hvxKEz9lO6zQITg5aIXSHSp+F0mraBuFEWH+aUPQ2vcTzVYjpD
8cp9zG8L7vfXVyYUx2bq1hw8QaSq2MW7Rso4S0OPFSvil1RRasjPi8EIe2DPPpVyrcrciWFLUJxZ
FFxqOhosOQHsNBknnbAMt7Z0UJ4xNv4/r5GRpow8Xq+TWUs/Bvq0pCEfNQpSMbxGwvjRHewrojAs
BlJyyf43Zk3Fwur4IMF73nxSpZxu+nBy587NuUw0ZDQleSkETThuUVdRFJkSVtQx2QSCsZYF4mPw
Lf40wWs08vtEY6airuK7r+MunKgiZok9sSOE0+IA3IMjBPscm+lVpf9+NrOD9dmGxUgZbrUuRGU4
gYODiYXS3IxBAZM2WjiPnNJXdbpveM3bsWsN0M8Gx/AvukOkgmQao0DTHjgQ9KWekGr1PBox9rZb
V4XTETUf5D0HR7XJoCsxAHx/rTEeTfKdPut8oNH/izIm25fHpz9GtoNvB+GvaIj1gapNDnKnZ7so
a/IlqIJeHYx7EGVhZLDdMvAYfBDvBWIsnt1NJZAOD8zDz7qouEULik/k3YIy4C3FAN/kgaD27/68
pyr4vJGodm/oJBLrICh706OdYmc4+4mk6d3EPiYzakv+rY2lIjGsBBifwx3rQ1H6aT3q69KK7yd0
YpTVIAACLMQxv+D31Srgs4awxqQRgBuZ8pfRKRjURKn18BEaFv4uwvBCUohdBt5WruevdXpX+7Sa
dvuO/qKh5oRK8inSnGcCL41UidyXaRzjurhcQdJIscZlR+xjHu+aFtb0NA/Kjiq7lo5khyTPmXOX
74xZIJD5JABqFkB+SloobhQMeJtU4tn2kyRT+Fyis5ujwCE5NtlzzKG/Ozi/mWfb3X4XPl/8lrvD
0eOnFKapCk7B5O9TiSYUv+/viEEXZ6pN0gtBJv1uodUsbBxtfzgNzY7UA2fW/ZjiTEvkwBlgTrM=
`protect end_protected
