-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
d+/PteVLKhvokt0RE+X/YG44gZdxlBH96VqZ02rSxVHgxCHAeNst9qAWsIjNsLAv5klD9J76xM3m
4VkAfgXYarSjemZU2kBwAjggk12cLBv4nkRqEyA8RA/CeouXa7ITx3rAe/1mldS2BVEEQwkoQVTH
YWLfvB9LkhZQTFxPOkD7i34yUYjPN7pydC9bIhpRaMdORhRj5lnmsDHLachmCvRcYZSF/yS6Q3PE
D5hwUSsUwg/kYUaQht14hkyINK3T4sbQxmeg44TApbOYDM/WYLC9NzOBXXukk97bi52G1w0Xi0M4
PSFxjJE9EWuz6X1UjKQ0C0IA2ErZx5WmMeT7xw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 17024)
`protect data_block
+M3/Jnqb/FRW6ZtChTKhYbsl4rPmexfa8r0dezS+qQzWVmnir7Tp+/eEzxcvGL2LEYhkjy85kFiI
MrYPXLAVYL5j7avVOQMOBRHMuDgh8GBctl6jiUYoigMD3VIBqMnZ9Lm1SjbjZE4mZAzn1CkQvPNM
8JNaNeBlp6UpjfE1r0fdoA/6aRDGSylic6I9iIK6q3k9zOqt/uaZhBZaSilnMCUROZWBo5XmmMo6
MAgmTvcOaZsaAEMqogENtMXFWXnfttwk0PqkDw9ibYtXDQn2KRoSP0fDAzGWSX9nqZW1zlypWSz6
TK5FyZ4Z8TLVtBo1GejZgqs/JbP8emQ8jL/boQua/m2/x1PCYDw0wUdWNLXIikGB7HahKJ9xFOgV
u63hz/HIXV4v8oK+W4NYJobIBDXndPxAUqv5Sj07DrNbLutrvmvLwD2juJrEXDfs2aQ+0VgBC+q3
pOhazPxOA/LEi7xrJf4cEPGcBPuMwqknO0mqFGL2C6sv8PTKkk8HjrqrUFSUG6W4TmWOUkoJ3E3d
j0C1/DZsJ/4tU7n/WFhiZFHoRfkoBGO7U18GJEyEG//HHmOfxX9SXAfV2R41hBfZbaPqS+4bvrQ+
w+PAB98b9UGqCanTOnDMCioGWlKMQeoD4N/Xe31gD3rLe2mWn8tCWSNaJTs7yHQjQnLMwrCafiyz
a8TYOpeL0dwfUk/ixXfgsDHbkzQjU50RX+ygE9huLUmUgjL6+Vui4PL5jH9CcRcO5o5of1tR7km2
iep2sEQlU+Upk6kGGxazPFMg7edsslf8whXUZQo/ycK5PpWDbBklQz8zIFpex+/qQ/UAuxr9B2Qn
r+192x+24Ku40n8DVuoiAytyUi0sPRIAxdRIzBnjNtuAL6gwaPP4ava7UJXR5zZYsx1nwGFuRVTt
DLR2BtDPZVzdjusUtU4rv3X+VvN8OPWtD4LLgL+Wmk4CNxLIfWnrUkXZjLRCqIdl2bz0IvTSUHkN
8IFmKLT2E/2EISgxrRRF8M8edbBcBO1etw1Mlzw7RAZtGMfkOxGCsMy0BFceX2nEiZqGfeD87yww
Nz1fEXoiN3PjDkV+t1Eq9oAHPD0oZAZqWl0OtvJLN1YuhruxyDp4OT7m+Icgog4Gm4Nnb1l1n+jk
uDgBOIv45NgLhUS6ZzafnNTvgIp466/A5IuUEWnpoK4kCBrdVJ/eXkaJ6pg/VSUOUY8FgMIjgqZg
yI4QCrH9aiAQ/ONvmj/aIVV1hxVE4CmgGG0OTEGhFFps4wt8ScKBE/G0a9fbmRgXDsjAu6/QNDD2
ftQ85uOQbEGZ4jeJkaljqBzMX/Vi4ogi5o6bVzNU2iWAzILE2wHzvwHpstLKZRY5VVnoA+7uFIJ5
gitSqi4M3cPk2NnMvwGkl64RUeCX7QM58/7qkct9tpyOCNREaqKYIE39cEqOGwI5aspGMOhsyDgv
ui4NBtt+HjYzH+7ySJMsRMeqtYmxapOZC4l/UHSNbR4FcmU7sxrYMr+oRstOvpVlPyv4NcFfguN2
aVoykPqg7oIgoaOojMUKIosCYKo71FFoQHG5rzLDXvwi7BlAe6Yks9XKMhIxbNGL8bhjKDL9iRF0
2YvO0gWIAtOP8t91dYGeknmcNY7jVajtMBEHU0xcRcdz+pzxNFcJe47K1iW7rh6O+SEMMGY+KDyi
5W0NrlyttOWdZxTR/USxYcvb0hZL8ie92X+qlZ43pfnb1on3/SDduo98aiNBDVDcfhe+cqkr8LTz
I/FqHxmCog6/CsUIGv7V4F0cOU7dA6kXkMGl9vgIwToPocz4R2Gtitr1VJreyefy26whs5gp+elS
PpI0FyItQoC/9RcO1mdBlsCgsSkX3YXh0ks/uTQDeQVM+dSfKGvPp7ok0mbt6fILi+XznlOn8XBs
+O7qL2ZdMx8I5jXGEcGrwTQKzpbyrH2rqhBqrOlGSqbOHsPAEvfcryukgrH+RAgpDPuiFHh1ftFP
tBUE9YOD4QNgoaf22dLxck/lbt4FADCCJUQdJ7u155NksHQnIL1TkLENxpOP6GFrq2a28+34o6HX
fL4Cvz6vM/n0r7KjakIChPWDUlHK3GFHCP6PcsPJCrBIWS7YAg7OJD34RWX3DHwCUxvsxu8esi9m
PVQMBfP1Mk9m0sDU8HK9OUtNhTX4yfa1MiB4NkWW6K3nDYNd/oNDkfuIq/T4KDanMLLhIhfwM/+i
2FyfCYeT21k6kXHuaWy5oyNQdz5Db2Igd1AcSFHNEUTd549mIVOMMYlz3JBRjgjU0FZsZTKs15ex
WInddBwHZcEOuSvIGImQiyqXgSlQj8Ox6i5Vmrfz5VxhfIeKLDoVrwTMkIlGfKTb0yOaI6M4q8wH
HQWcvxBv6BbbjVQCy15laCuW5H/vGikfExl7L4UOVG26+ervqOg1dU2p3qJBSZHnWN3Dzh5NpBlC
0tzLVUogCLIYq81nblmeFl67G+Rg9r+Oww23/ArfnDYTcw+95MawN1ThUR6/z96dKZEGaPVXCXaI
ubZXp9Nw/9vC81R8uqekLObCOrrnMECdpGLIMtM3nYEudTItLvivAfrrLT8nu47I+K03PbNxf+Gk
AoU8omIrotGo28xsCWPj7MnJqcAqEI/Zq19/ztrI9EMgSzAhhyIhy8gg+wbcrGw4K4TLeoLwwz8p
GPJCscrFFCxu83M63oRfCyLDfeoqtFPTepxH/3J05esAUqVQti5kTKkA3k3IeBNylLglogR49l/Y
/ExWCXzAqcnzgQuSRopCnEPimsawJmFM8+gHPSZ3hAJ/l1II3cMmteYioBqG1KE8JQhhAdCPLEsi
cpuogTq4wGF44VYLyeMVj3Ei6h5knfOR63ig+rlplFBkrregrO5tT4L0m6dvhSw9q+Psb4hhK/3O
T+fswtdQZF5xdCtvsVddcPbmcxSzkoXJaEqrxM7TaBOuNDccEQZrzEnEaTGyuHpy4jfvENA6P9CA
Q1PttSVENq8z8kfm9xf1nZ2bk+msZOJBUPhcPrsPY1GU+b7OtoAztIrr3twV3+4GbyVghplVrH5e
jjyhlCSPr3cyF+eoFJrwkLxlcJggWoL7LOI+cIMypricwWZvd2rwrHeZZDn+LyJb4FReNfGD6WZc
QPs9mc0ftTEXQdCXurEspbu13bBPFDl8EOI8wBlQJFtVGNNmfpjQTuCNc1j0iluAfeRXy+rdixgq
PP308/fdzx0+2GOE8tLKXub8SmEPFnnFqvCwdEUMoZTnLWpQZMdNvYwgMCvVKrqMDEqteeMFC6/u
87Wxe7KFwUc+iUF63datQSoA+4JVQCphUIZjohK6UL5vfjzf7XKZN/ORgpxoELzvTouJ/ckyxqG/
1nlYNF1rL1oah+5xgUn/Jr5WIy1MyVLea7i695SC0xUfFQgAa0sar0XHUpgROQRhCRIvBPISj4B0
y7iQS1FkAQm/PkKU46rsHR0KHRlzemcDEaZH7gRjF5ZRLmKctFUcWWzHuwgMS0m/BACFwqUS8Qsw
H1DH5ePlyeBsr5zW2mgLVvPgBiKxYoQdfyc0sCLycJk2ZFoTOKyZk0hctYFEy7M6BwUJRbXDumXC
iSluZMEYfdyGHUqleDmoYhsh+juuAsC8oOGEyZabCbRKoaewRaxLieKQ6zUyneiuysSqc9b9YTFj
AHIwErl0uxRTWQwD4rhBuPzZpn6Ez9hsmETs+9sL9jseofik1kYP7iTylTRXSVL8jEEuAm1j0DgZ
g0woDPey6yGrIjBN0k/cAzDbaU7bGk6wOs1Me29AexQOL0obKaYzBpUW+FbKo6ppezF0rCSaSTkD
S0omqKzvBESaJ0ZWTYOwMsy4C192MHol5y6gVfoARZBla5QAFWTQSA+xmGPpGbaA/k8EU0oPbN/X
YEv8jS18Jy2aNkq9N79lOZ2Bgb4N5IEh5c1AvTPpVAKLt0FAZEq1kSrumc/Rsu+SSMm8zQ36DgfO
3pTN31UOTDQw9/th/vIaPKcGo3c+jH9aCWlk8xv13Ucb+9RsQW1KGSsJVZ3+O2EBfJgw/esuPZOJ
pZBZoQakRF9ddF6shYTJpU2BEsH1Tfj9m8YbrHo+nn70MJiatkg+w51XdBr7EHZuISBdCBlmqVaW
vfxWPArWbEUTXPjYCqeICQogstMpm7eMWTIVtNUjMY9RxX4DHAbAgtUpljMpRnukPESe/eYnhxaa
tNxjrih4/nfB9P7hDkLEORnXty7T7eB0ZTi+TBMGikCcWIWjWSsnqAC2xJ3Wbfif0cIbrssujL08
bMS/sR2KUlw0j8fbDUwrtnpqdmAEHtFP5on8CAfNEEOHeOK3TWRTl5uFO+3P9l9JNDOcGO+0qTp8
Fpb5KPqYLGPkSAbYYtx1ZG4HHYsFR3qWBGr7uab7d9uigh4rG31cEGvfXDJCk0M8PWMXqsg0nmpc
l7mI+J7qnti0RN9Oa4fsFGBh9PVdWH0erPSC5RrPsjqAatT3MH4bCCWGeerKo5R4x30a6MqgR6R1
1Rs483fve2CZ4MuqOfIc/vjt1qzdVbHcE28OfFmyB8MMFcizBcZdDy9gQqz3KSPmzO8wavJH0ETc
YWbyKkenFL7JF99re2b954EO6JuYFLT9DsmX0kb/nibQ+krcUr+gR6gGbrNpE6jG0sV4Wefmw6h+
RsckhZbSHaJc0mx+i7omrvZHKkkXhcBMQpYkRbk+FoZ0XaAcEB0/TER7fJDKqimVCBDbE4YP2fZw
oqx9+HNUHXBc/J9Hg39VbW36PyuMazF2QG6ytFFJGA9EPtSrPBGYOSTMeSakBZvC+fABlLd0uRXq
TDWUnyoebuL4lUiGNxqc7oEQJ35/vrsp+5sNdzPACXn713ohUtHIHoGsZlnq0zIUAwje1lvTizk4
UH/pzhVnf7NInbbHQ6OncxCz9e7jbkmCAmTpXPEjOChQbkGmsidknnsGcLEovcJx4OAPOMTFOT3f
qVSSUdi2cOc82//7YepyPAghrRCrSThhSqHqZP2e+OqPZrDzevyME8uNDL9mRJxnSWwZBMyddWXz
9oYQMsjzHAhQEiFDSpsSIFRg+8lvoOB1vPSQfRPV/4GT9hA+dhIQ5v/PQl018q8Vl8t1WRwGS7/F
9zn2YRwaekljPy38BjADbrfGyh0JR4Ju2R4Nq1c/PK36DufgvNzDJakaELC6NAkTCdV+sRtbO88P
6dIqb80NnxLv8Z3FbY5qNtKA+7I9Qy9ZJeBQTWpPWMIQJ9Q6YXOipBn5iHsqWcN4H2GwT5Nu4maZ
bM/cUSdp7AT4IRuLCnLD0ISktEpNdOGVKDNZesO+duAFeP/xzgaoy1QXk2ydqxnaJRpHWHr3PpQJ
i8o1Qv8ietZeaBGhldkY6pCWEHeeQuq+bdz1W5oKbLwwK4n8H2ibeNhWTn1pwtCm9jtRRqK/jLbB
DGPzaAfPt2rmVqTe6+KuycPRP89QnIDw4PHFO4vl7/NaGuFwO9295nQ+xkuVSUIGTo2JcoSaqLdz
GVk332ybxazmG5qgOAIR/LIL85XkAC97JDcKLDRPlKTyMoiuwvMedsio0yAUU9vMEQzKWGjO/rn6
XP6nDuq1NIDnwPbyBumR1KDssaaqwS57j0Qel9Nlw6WPTEyXhnNy5GxpcZVnedLjQyoYoPgcS4wI
uYAw+U5mynMwrucNuMa8To0klJGZOollpBS4AiNuXDM5EvXtwfmorzikXUNTZ+pCjc9kL503QQIF
XhOcEE4fqY3WjzwfXfnKnzEGN9ctn44MQY8A8p3QC7PKH4wEtGlfx+1e/v09pYlsdugFzJfyQI//
Rx9N1HYqKUhhvaqnQ1ky3po2XPp7+b53+QUlKHSZH9i+DRUbPKDVAX2ADtR0zZ/WW4RJOFotSTMe
7d0A4QBA2oLrm8SrCau716I5l2nx8+eg8YtCyyHodYRxot7S2iHoV0SOKQD+s18EnleO87L2CbtY
Y29tUZswRx3FZE161MzowoCZXihbW4l4E+DJraG7VZtY+e6lM+IFhsQUoxwS5pO0CdMPhkwPkHHT
A9+0qcJ2l3QaA01Vs6lkM7wBahLhtoOD8fOuzDULCe7hsLImc5k3BGcmxjvxLvYCUVtPTWwquZzE
pzPtzOdtUsLjh9EpB/dvIuEqkhS2vJswuMMLs3b09xucPy6KHvlnOzFeySR+5rEinGmLKe8oSmU0
PaNqx28Y2sjaI7WkgG45zp8NhCQNMxKJJMJK+2V3l+ZczSfS+j/BW5+fnx/fDcc9tgDl9hXGrZnh
fFY9CSkA+yiDNx6fKR4k1bZL1BTzeZRVlW2M7pMTUvtJn5AvF+9Bpfh6DlVgp49MRmmTC9gi3Inh
eoIffnn26FhkKTAH5FD+W0QCuXzZ9jX1iHC9SbJWEJ42WxWo5DIFatjQNNDvsI4H5E/jOvkX2s2N
i4rjUQieeqEuKWvxEpRucof3r0ih1I6KeTPwns+1sMAidBJ6gYA2nghRu7IHUCPO10n3Rteo7kUp
EwEKuQWnuu5y2GEXHA6e38CHUUYlTQlZY23Uaqbh5RvYHPGReND23gfjw/pvCONcwI6OuMvl02rg
GnRPQaayp32cJIIYriiCDeuzC+ys0SqVY06kGFnsqgmpOVIZpXdXmRZXnO6ZNbZKc9GdWNw41721
rb7BSyvK/N/9l+duv7uLq3E/w20QLz7nS+zDtTpafyRWch6YdJbx5hik7wqq7gTKU7jEEfOxCzEs
yMumTFe7iCw7vDMzGUVZ4R1E2CyLMXPZBCjTDx0c7NwBZafMTD6MzpQx3DI0FnjHsMmyophE0ygU
sL8ItqYTZkYZLmibNTLqstgxnkpwk6K3spF43PJQDcqL3wthb+XWJen2bap0KgAfMG1+e4ybkBcS
/KntRSBnaW9GbTWgLo+IF5OMwlxMX6khlHe+MKTGUVIiPbzJkUTXIWB6zh3GXonnX2U3Dus60u1C
4W9nBod9ijgkYU55cevehi0ZuRcRye4E2MlPpaGUragvW6361hoamWbjt3hbvObqGg8M8vYYpB0f
Q7qLlJl4ONOaxOLNpWg0V2RzJHzqokIZs1h+1v22ZUPoT0JgZrYtQJJnRMXZ7TJXdCMjPDbhncbJ
W+9n9YBEsy3o8JV3dA0yFVYEjRHr18KML6N16m7z7/qbqin7f9puxm2Kw8Rhc0oJhWsU/tmTBiGT
8GLEjwtCht867Bq/POm6+bkbZAfN6J2CkhRJHmUl1U/yllJi+LkAX8/J+BovGFie8kktSwYjZlDF
7F8GAXSipgXlC8gDkBZwRNTF5vW4PPozjqnd9b5kYr2DqsNu/ykWuSOPJUpdKHOm/x6VXS5SyUfL
elk8Dd34zUP2J8HvcueChBjZYP4Gfv+AKR2rR4y1IN/Rv7WVwSmrAqy58jh+V0G3vDxm+Zv+HRV5
Puyye0vNF1EfJQpRt+3XlAu6C8EW7hh4Yavw0+JJI6SqbsmFDkuDAZdtGExhQqMDe26lQCMed2Oy
+6qXaDf2HpQk2f/zk/QW9r08eFppoRATkUr6tfBkTRGOujPDamVng1uqwPjinB4Z4m9vapcS3yAA
STY535PoDQqMO6aVKQzWNKN+XVpP5UzkRrnz73WH5W+zb5bN3RlX22eBOF6FXoemRrIt2mAcWt5x
P6IRLsp61Eq/5cxv2ZwDAY/QrvZi5Ncp52BMaf9Q68XRF4o1R4eQfKSoUGFMHzXf8cBTgVjxJ+nw
BZM+FYI5yuY9/GW1MQWdw182ydO/qEDINFMBodnJCfp5DA+0ossJnQv7flVDkWstdRG0K1WXY90D
gT9GzEt87HiRgHNx0yZ7XsCrcz8HiALetTQyjJX/rOJZGvBgXWktUyHr9hAj/MZEP2WXpEj71lSP
cFeShrvXONE/Ip82bAmC+d/MrCmwv3pKZnIxgk4ezLbi7uOBImpUKwt0xZTgX9F8rsR4qmflTpRw
SpFB7kA4ivtN/SmRIAzeYyC2rA7VW8XlrdLPujdXmJI1TB+QTOH31yAW18Zn9Vi3t4+zD2kbnt0i
0Ry6KohljUif9LqDgSe+NGPc5hyTDJZ//U0eMLPs8Pqggve7wtm2ogsNv3p7MLWfgUk3968K6liO
9qnEI6PH/0WW4a0bcb+NoY1zotWqJ69uU+4Ovrk4eRbYp/fvUbvT+M2mVK20RJIDsdkuxCp1CgkW
BOldS5H5lORRjGPetq+aFnIXGbIoa9KZwWGIsucktLeoOsu1hMCPrONaqfC6YHMRKrnNozAyISzA
vayPv7e2p4jNksv75pUYh897LiIn1qVsgc/AIinwBMP2HWUSfsl2522rCwj/aaPYy9A12BAsu7kt
Ly5GMVxq+3BYCkwB0mBqO7ov0+AwdYtw5XwafypP+MHAOUcCOLk0REwY8lnZZhNc6ih16bMSWrpP
BZXxALlNjGsXl1eDShiHd0dNjQOnqA119hqYE3TSlvJlUHH4VTNyQ3QNaE2evZ6kCXzcIULFUvvO
LqWEnREu2FT86mpC3Vgwr+CVajMnveie/554AG81WifGSVcX5hIWaPJM/YAnkke5KE9tz56HtOqk
shZO4jbY9pqEwXrYe1wBVb98HRfuLCeeBR+IvwaXCUJFQC3K2UVgFNpcavrbQEUkmzBYg+Uy9iuW
4fOrQSdK4uEmdsMp6AQJhiYPow1HcCcFdcxQEPm0KlPfkALYQgfjazQrpJoqDBIBqYfXzHepnqXL
i898/N5jjgtFb+WmADO2FQc0HIO4NmFGldvZ3j+pSN7QkRnSPvUz4rJMsy0Q/SI60uK5WNaHF2Kz
CLyqmau8sE/rYPFoJiGKwAb3tecAl9vsebzZCkY3FqArZ8etdGHrdV6oROebEf+qQaoPnwG6aY4Z
WOjKFUM/j2l8u7AFF3mTYyKFqv5oUPn4MyZrt+GbCfvI4qVVU8u19AnsSo7viXf+BcUHqDEPFafr
oSbWra9xYEeunf4qNCD56Sput/8taiZvqWIT/YqnBKcEQkTuQh7mb0dunTzjK6P27d+ClZV5p1Wr
5ojLlRllLNtUY8XHgGAevOlaX1zqZ5+iAYLDA+Mc/SdoZZAXkZe0+//T8XPq2tkHUA0LphTO1hJS
MUuJqWhohFdV+r/0vs0lqBgLP3xJ8mbW7GdJIbGl+1+I8Z1d90ZVmobkmWEBA57C+jV/XhxzDCPI
xlavyQv3AXMm89pLPrXGo9T57hUKGRguElvo3W7++BXY7uhpo/VIf+dNc6LZgD7uPF6kS+p9+Jc3
buJTuH4MFM32Ui2XFPrsk5oMuKChgkvK1Dc7fkxUX8IDNvFDtDFsMV9o1jBxXZ5AyIkHgvu4bza3
rS7wLoeylq4csRtMzm44HwanyNA2y/WPLe0HFLxz42V8wLtByYHc2nQ5NrXBmEmrjsHiMs9OTrvW
DFVAD7XV15w4a46RNOAQ5WkwsWCZDv4IhPplxzEWox7pT7fyCjxxknDniCR1k3lpvdm3m0wN6Xw+
p+rr6WUpE9CJ43EG2jPDXjxEh7pGPXDpYwsPVsg5jmpKeoxc4ItTZj1T/Clg/tURl6brJd1TvqD3
0uwpGOcdo1Zcic9XaGqfy6MOK6n1txlGaXnvEoDrw5Z+3RsX7CFkLZZKtWJhh5BOuHxfK8eV92mh
FG7tTCPaDzIQy8hBtUgsEnG2iuuddTS5UzH5ZaKb+7iIK+WzLT8avkohw7znZrlT5raHw/B9EX0I
17OE/mVqi7AJA3MO+FBu8NYnQOTCkc5p85z4wNPHnfcFFQ2Z+WDOMfrpAr6uB35V5yLGUyt3lGBg
Tq98O/w7AwJlXrL771Yg/95fpA8WPoK6ZG7hfvfcNRSpzKG0zBSHf9OZMnKa46YNNK9wTDJlKDnk
tY4wTaF+yF8V9XDyxHCnRi+jVz6zCF2SYpSrDOabHQS58cTdgfDwN+M3icZ6TqfgOddg9F17RS1+
YUTMmtJYZwD5e50km1lif4MRP6sYpxZU1MUXW2Uo6jlGU/iZuHt8rXkS1ymj9e99G8JrNxAt4Obq
+F+vwOqoVVLdsBWgqjRl6yQY0JEwBzfmqv4tuVFtP25c8FV9MkcsEydUuKqqyO7owAFHwz1U4J9u
cbSBw+lnmklNimONkHniuXKOKGZCYPkoyssVQF1M2uGI3R9DCzTBv96ZqUXgnjmSosPH9h89Idpx
/aL7PVUGXrplLIU38KRlLtbeGXU8dPeT4xyAnaOJYnA08vsdixsCyXHrYH0QH2dZSG4DoNAVnyc0
oPU99/TkVAMkKNhuEhweATAEPq1JJw8WiAvLZkfnASM1fxt4hGNiHvCTMIAeLf22VAhKmK+ckbUS
GZI85plc9U6u0TBvalp0I66PAqeRXoGRr5wJeF8E7SAi/cyBLnkexUWUUihhNRepvR4ksqEbQNQ2
P2KN3AxNSE8DkXu6tCcSbkpFOV2j8CVrqI35Qt3vRQhrGDOTy77h8P8mBvqDX/NIStV9OdR1NQre
Tf5qc33fiK7ZTFUEfMbHouqZIp10lzNhKaDvpJNrZCWs9tc6SqsXXfnIKOxbTFBoz0SYKjyaCHcC
IRPzbCNyI0aAti+W/TMUPJtCTkvEzw0YsSDVwiXVJyZrzM5YbQhVYP97zMD9oj/0rtud6oTpE3KQ
CwO3WSjFLZlVQgjYj9RVuoCyFdN9bza7uRCx34AyZKyfiIOffX7dkWCerXegBjw3IT2F7yV7GfCV
QeKfTRHM+tOhZPxc1gmm7gBZYugvnjLWfOkev9aMFFuZzvqa0dTYxr9h10qqkfjumXguvqHuG80Z
SEAoAcpkCDPOGuCvcvP9sQTWe1NMxLgX7ZC6QAA/kuGfgaKO7mYiYH/ME2J7oVjwf6IfDXWUg3Er
lzOnDtz2k9xPq7auWgB7imGMSQ6f3+b+lBI4Pm/sz9WM4Ql3c/FzpnWU7Q9PgrxpYYrgxTb5HBGp
BMiOcCvaW9PwxFUcV45Kg4IdL6b3Gr5wQwHNmN2cOI0uU9LmIlTXbYHwcn/qYXRreAKX9tnoZKIl
8bK7f9hZ196Li1blbb4XTcK2R9OITminPb81b20UmBgnbHF4V2qAlsM/IDMsahd53q4JugrI1KIb
BJCBdoRqwHVkUJEHokRUmM4HCd3n6m+3ym9e4IqDii5Jnuv6t4za7Hq1WgQYI0RydxFyyq8V6k1e
10Pz1NmSCvV9OWMtq8m8KKWWtp0Fm/0uqX1SXFXhQy2Ibg4cSSLnzlUG5bAVZDO1fwFSeiVsh7YJ
pTMI1j1GSgieDBHrRaaOQq4z+emboFXF8m4cbWEaJ5ZB6MbKWy8rzffT30U9U91IuyOGKv1GgIqG
1XPfPRGa0myVWMEG+EbFp76hTnFR7sIxiZbRef0p9lFpGQgBSm98ZIEjqUI7Oj1pbam2ejlCtzyf
d5a/ZxhQldiRKVZ0IfjPMZR6YcZTiG99G5eK8Cgf3d/syBpJsm/e6W3FUqvN9s5fEb/x1JAuLXPE
Ln2a3DWnmn8N+FYoLINOHHmNoj9wIoqVKjpXm32G7c2WNBBIhzmYMJDGVh6yafGtBAhgIhVlR3XF
F9RcwSELtz4P6HardppkMbvUvZ3Ho+YkKfUEbxDy/UghTK/zstFXqNjL2VukHdceDy8fqmk37C2W
IQQNphgVMgfxJQZG67/C4zn31aFpYqLYu1xiH0wuvrg/ZkuLWn8z+taVjYAyLddw1zazh2ScVGag
WbIC5wmtv1hTYqbFRUuo/9kJNgkHbSjZOzGf1Tj2d3tdsLvhC2xAQOWlhk0LUter1qM7UQhYdqRO
+C+cmaxc8v2SGjyO90rHQNskSsshReg/bIi8Gsy+qQXCy464L4CUxC71nsQNBK2zbFDt/P+YpOdz
Sbvh8oYaZnOIhUl1YH7QZIg04lLkuX7uRoq+gLG8UIT4MqsSaSo8jp2PM3OSKDCeQCslrc7h8RfT
FZedN5BEhLpnUZt2cuHeaC6msnO8FKdqZX4clLnt75Vh1fapWTfi4XCmvezrQt+m3GR2SCuKg6Wr
B0LdF9KsBNZXVYFXfvNDDTWW+E9a8Od2DMymgbXRArtBHc8I00pCYSIJDOzGoMjdNzxanNWi/kjK
nQ3FBC+R4CR1ZJ5Tpmw5asrKn7kMGKOux21WCWie0rL+acU99CkZkuzHmwrSfx5e3hJ8/I7/DWSo
ZjfnfN1ywKDT+yBdgom+hONsl6ulUShJgSQvqKT6L4pAkCySTYUTP7uWJY04ohMizR2NwBIwC2mY
pWJrVuZij5y+OQSYhIIX3uVS3Z4B/uxcJl0skS4/BDaG/JBaLeDhwfFojHjQWjH0X6YHdM233zvS
rbCLOrNrJrLVarGOuBMIZrQc2+sgtElgQXAU+EtwtFuuBTVi9CIf9ZVJuWbcMHtT1JykSl3gzOOm
Y9UQstg+tDLg7xDHSg7ClyPMzhWjD+7Gm5FSzV0q05pZ3XdIIwv35j0TDULB80aP/4YGRCE/67GO
muxIK278KypnDdOGp2kJubMS0JWf5tRQV+IvtR59XSG+dEfSX/wbTOHIt+aR57MUNqkgiI7G64QD
6+jzxEJZ8OdxR/WbVH+AaFRiDit/scnGuJBgq2MU3W8AzlihENV6nddcSjntkduAmpYLHL7kTmRF
TKe7LCPTDZ07sEaLg1efMxNtrvNESKgCCv5QeCfAkRXbZdtKlLlRZBp+nSRUwcuLLXtcNFo6vq02
j3uyNyw6irb/mCKe9Ttn//UABW9WsSMw8zEjZ0FKsTztuIOTLLstMKJK0eyDVp61pzE43BxGylty
q/qX/CMYNV3yj3BdmQs3HMhysLqbsEu7+r1MiWoIHmtidItJDYnZGHoTRAoLRuZxOT3iXVWy4Bzv
iShx/l1d5h0BssYS3n/ju4qI6bcHGsjWmVu4yQmHUbo5h1R8xF5RZ4EisWi73rZ02gj2sLwJ017q
hpKL2wl5T0+tqy838Gpxzdf1qv9CepYIZBQoRXGPNVUtX8hXqGsThOlrWA2W6BuiK0lW0rrOhc9B
S8z6tJ4rI7d/Zbip28zUMCKdTWBf0cF3ubD3yRiDG4fLpQCjN9Q05a+qxQhlPb/WkL0cqI31hNlP
lWTZApK7Ubj8Q3rkp99DU09v9k8GK7ySuxrF43j8TgY3u7r+vU8YuTzHdhoJXUQ3/V5vXSGNGlTm
biPX0riU0+6FlVRj0NOn9jQ+vVaUN5JP9kgGAM3vTEjY2mYdU7gB+0Pj1krOfOBus5IhBbWfQcgZ
PAAap8Gm5j6hssFyNKtK6QHCe9xtMEJHGuxk5J8zYNlAa/vd9XOtKe2EUlzWxW5Rfcfs+ZlCGMsC
t6l4E7pN8hXET/uOQu7voCn8sN6p7v05YHs1uV5Majx8hMLFGRwKI375SOyi9k/BHhFHdfFuHQ50
FeaCYkRCzpmCN5Gn5bgTPFa313EV7TyOWiG44Wv3y+lHh+XYepdeSwdspzKLQvkyAcySLy/DPZOd
4CpUbh4m2wwKyfM5z3JsEUVEqg6wjFwQIrnsqOSApKkplQTImQeDIaOICC2yOhjrLL2dACAoYcbw
DVMKyK/IFy6p9dZKTXDS9F4KSL+msCTdSLqimHV9kjpwEkCCgY+bQ9LZQvmJUsIxi0WG5Y9K+RW9
l3fuIHZpHbzfWPbrCVAdl2WGPkI4RhpS2uUvzDfv3wSaT5OwdgtvONojfCED3SrwOIZzGWPDEckH
69tMB62EzNvj1acteSY9dRwdnGCtxwVjvC8JoQw+ohkaj7P5CmtAtyzoCRVemBpdaO/wC0JZgZQD
BQRVBH4zskBRl/DbmQJzY33A2vyABESzTBj0HwGsy5wRrfTX9g/D6udsADHIUyIvmbgVHWOfLo23
RR2pm8K3y77rFhP5zyr9YEDGXqEubuSMXV69Hc7vpCV67+/I2C7QYbi9DTAK37ShuDi0sjJQSowO
uIPml/ZdcDfTa220bdz0dScBR7+rTIgT5e+RPt6zRL0+B8F7bAWmfkknUfqVyxwxx++pRUrq7FIx
I6SgRvXEM1WO9mGBijOJUfx81Wmc05klkK52O7a8lhSD1PhBheUkOLTdIVWmxOD6XvzRfcCOjlMU
h3LqrqOKlYGA1x2K1SbMspwGiEaYCOJFVJ93YuXlwYXSvpm10PZwE1MRjCQnCRfxfVlD5aKKEiQU
ucYTp3d7LNFwrVhMXoNWODns1pPbTDNgSfXzFmBcswrRQBpQoGHdfXAuqzbfIzYDO+DZ3EOkyu9u
tb0C6syPbVrBodOdxbuSDfV117oS8dkkjRziNnkVJxP3DoNZuL/A//CG7+Ch1tQUObvyJ8hR2R8S
IGUsx9f0KObNMZmJ8ASb+1GYKfhXr597KVd+6+QpoMyY89ZSAygno2k/9NCkP3Wov3GkahtRXovd
OAMLQggkBhlb8UFRhaKMvu7+nPOZxf0fDx+r6Ywq76L70tqin1uPvR7xcfvWXyiJWduFRUPmuw5D
kHb7gDInMYPTo5jCL5N7LuPMQJkbi0SLHQ24lzKvOhjfQaYPB02/3KmkTqXLWukYiAQE4dS0UEU4
IIP1Rxc2UIYVzNkfKEkMd5bnVFZJpOG995N7wpshQMhxu9t54+FoHLbx5ROAxvQO65pbEtZnRpbe
oGjxQOYflp3Ktv1wLSQ9CEh6CD0ItpJQGI3E1DtTDP+3DwxKmLJlMaEQGDHXufMte6/AnnGwZaXH
2BxfkXrsWOhnvm5CqEn07SulcrM5gXnoplSrGckw5jOHRhCgSL/ibO/CShb2Ly9iYjZ15bL5Ml1A
xtD81JLOZqrPvyAoJBfmJv/5uHtXpsBA6NRv4XwxkS5WrKQGwQSwgu1hGGnUxgD3E1lRcz2pc5GL
1YunfOEgSBZ/GWiLKE24sTo2MBCBKPPXKg52XZbVNkGQw7t6ss9i3cD4UTM/JXbkTI01KP/ajb/4
yHfSlKBNIoEs4Gvv3I8SoVNu+B/1YLyL8my4q6io1Q0PQf5rx9wK3JOXVyjwwnOOpcdEWBt40jQ+
6vGLbZ8lN0Taq58mtjC0MGpVhaxY3UdzAsx2CeVqT5E/PSi8FqVP3ot0qRSniTuFCP1rcti4Mj0V
qdLiorOdwM+grdEqX3wJtEfAbb1m2oNBGwmyjIylmD6F2E6RNtLi8CqgdaOP6Q+UgHsQc0NQWrvi
mJsWyYDQxiugLo2a6OgEizk6RGr8y2wK81KYEHhIpA0trL6HZphnEMlAy1/94AOkGMvl2GnQWnVT
3wKVHkP0nPy76Sl+fwtE1m0fXcSjRKZZjpL+OEVNtOE0I2m709f7aBL9BH97lB4hlXHhICt/7GEG
kCXVTx8TJfBAgCj5DvU/YAXtlJHfKjQu6vLgmX87xzMfwdbjzoVz6G4T6F/xqVh+dWqbI4FY1Qbx
TVxtiq2vOWUzjioK6oODdL1s347EFhKyX98QDuO2YjSYNvwVcelCanhU6aI4cvM55grQsa735jWw
hPlkIS0txbs78Icb/5OwGfk1vXhwNRugZrEBVp1SdRdtJAf2RqteCZCROnibc+KN23j0uUsXiG/n
DPNXeYqq+0Gd6rUO5JHE484Gh6l7EvTw3Ad/SYXh8D0I2qJ3KlRaVQQ9EyP4wSm2iU6DbWg0W6Up
BHtmDY95aQbrap5tCVjn88H9DSTKPzxP0WzGWjrMIv+59JrM9QNLwDKF1ywsn3sbHg54x3tnQ+t7
30c/LWBDaN7uUKgGRzFDJuKetl1sjCD8eaKa5Vc1o+L+SkutkfcoJKszU3WI+mn3yeQ3cONDpnmY
wYHmE0XWdPcRKOhoN+B9IU7KciEpX1epA7ego8Pqh7mBAuZYRDRgSTnfNnCO1N0S0adEgqTVFXGR
VseXh/Ij95+qWdFbzM6bT5Ay+0H37iFnY+Nr9WaAMhse7SleR1/u0OdbLE0qZCylPoroT5NXNxJa
6ovKQaFphsmnIh272CoRw1cNoEmI6fYx0/zkYfCDzs6semBx7DJALKZCRJOVTHNtGmxwRf1tyVi9
y4Xd7/VQ4PUklwZPQUqAx1CNDbSFsrrGR0TO/cYKUrBqqGnAimOp4SqmDH0T8aA6x3/Q4pUmLoBd
28IndJgtych6pMmyaMjZEs2YNkYYXLqqYzFmhU3pJCkGSiOkCSTN0F/lGkHlLjyzyN4w/yT4kS4Y
3Z0I4Vmx1CCcAT9fjtLruOm59T75HatL2B/8eU7Ff0v50LgZlEwLimsr2g4iLJ/8IFpULKLEeH8S
zfOseur3QwXuGrZEBZL1ZIWKx1yRFlbk7YpKrPo5MhNkElRwJ3ALdYZ+3ssi4SZh5zP+SvMZeCEf
lf0LRcmSBpZXEyoKxxY4oF5T455x0Bh8TIBck7daIz2P1rMWwtc5uc//JGJzk3uGvdRMPlPsnDoR
eZNavedpxhDxWcR/WOaRNdnNLt6TJ3lmPuhNiwmhytwfYbu71B1fMhnp7jalghQhxVgut01XoJeo
NP+r5GM2yj3zLOBR1uSUcSxB6Asj2HReX7xNnvF3FCPNFAMOEYulf5zj9OgIYi/IWxnA+/eYuDvU
7zy/PPkF18L8kzGYyo0V8HpLNbtML/HdE+jhVmnI5diHCZaHXjCU8pGDFny4gByjsW4uCIK8qrZq
kRblL2RqEfqQUWVaFImQLV4J90GJrHnH6qV44bOo3FfbdxI6EIgslFDNAebYwnHZTtANp3UHjnX2
TJHE5QryQIQfxhuRYgl309nLwukbmxk9QVJDYt/PpkrW60dv4xU9sXIYSuQBiVObdg3Rh/VvRr47
1jGUVAgJiKwguwWz1xs9ugHU1+8kJeHG7wcd/uGFVdUiU3yDwdjwfvlv7vIoLUpnYhzis6USAHpx
R74KUanJ8U3CfSvg2FIC0mL5+9W/Ghkfu/pwYR/bursnpSxrDX5/vzPnzjsKe9NStdPABPt1+Rzn
CNYRP4sr3+80i+MYYKdmGxo0ru9z3j1ov7vrd04f2NJaWWHFqr5TzX7ywkg6QImwElLR/nBGPRoP
vNV9Rk8rt7KjMU/6CHrrBgdL5rGO6Za1u6dIPcJQRqs8aqSq3NIPgeD4qZ58G+ybF/qv3yM9IZr9
z1/EZBpJX0e6nwgAPkXBeAbV4QaUE1DD+bpqZ2nsn7PMiiHKfM/tbPdCTUoHAWS2LbYZP4/jPK2z
nYIFPTjbXm6SanfDbxj3IyzFYNH+GJKCmxLJIH20S6+f/bLGDlwGL6zXeUCzDa2GmxSnDbTFrJca
L4bVM7Bh4O40mhnE+RbFvetKk3q8mXI/2Yi8TMBHaTB1yMYnGSwoYivhlozrEJLo+KnejepcKCPc
LGepP2GU3Q8Hma96bBgnhWZxns3ruJs1+G6622cp3nE+84nxCHGzikV8lYUaibdt995aXAmBtRgZ
G1ro+B2V2596WgPSxYIg+4loMqSVUCip46Wqf8THk1ATPGDPt/pODS97t7+siidw8q6nNwEkKrI/
epJ3bX3o1krxjNCFTi0ZFAhcjEZBINvSn1lbpwkbdy7ORWhaHN54rQICkvHDK1d8MBGB6TJ7bNJY
VBZxkoixGhPqI0vQBGq1sLQRQlT0/l9n+kAYc7Q2rRZv7wwU27Xzy3+V/DPuPw1fuzDQcC75wlqQ
5J9awuVnOfzj4vZ0jhcOnj8BFw2LIdFwrc79ot/9b4M7qww4cfPoxnzSMr6Q6YJ/1OypQHYuRCrR
rn/xr58wJIGARyAek9wVNt+C2USJeXhTdVSzyu+37AqH7KqjnvK/JJaT2sMb1b2h5oiHZZlcnGvR
X8OPN03B4tnOfbDzxK5lwiHmmnCgkQUehJJpKfp+jagdmr3s5rRfRzVlwpYP/h0WlqVq1qTcitzq
V75s1W4l+JLgcp+qV7SHmLon3+/6ZYyPLVjCv1Lq4Se1R6uyfLB3whcOJkIN1DXHAR74DmI3+59y
49uFE0CILdjBhpHB018IA9V2p8KPmmwR3NmTdPBXm8cgofH6LRHkd0AW/Xam/94aqqek2xQo8wI/
MHIrA05NCce8uS5We+7h5w8QN9uGW4gQwG4Xpah7z4NsA2ekOfyj7HTX2xpenijUS/mkAnrmjBwY
Euq+AH80GtiVi3SOSdD1h0zzJN0gL5nwTLVFm2KiSh+zylW/4zdff8iOT/0YAEsyF7Dylg+tamPJ
Ozu2oq+LUGpc5w8x82QXEXN8G1xUdjwE4q4dJXjxTEdU1ZHbk/2qqumkrHgLqmJ5k61GI4CEbLDf
t1FC7fbpdGIOP/FU9CASBnWZEYBkbvTSas7QikEMyL1s2bHXlLgeHBROn86F/cpk8zf6kSFFGFDU
XpQOcYGUjLXtz2fAiCo5mORYvC8jupdcQ860iq800036mUZ4ATqmXzR6AMT4luXRLBVl/kVpSw4v
ZgWWI/GKpZCWt0VfBnl2ZkERRhZBc3YynFKilH7awCEN+ex3KQOtZKBBN6UEeUuhvsWY4ybYcm33
kQZrFifeBA18JMHzob4Q78Sd3g639t4sEj3g3JAHkgXdjUE9kLCssyFEYSlJO/n+Gw+5A9ebFeNz
E+UwK/IG4qrcnuChnygqPJxqdlBLNoId4252FcLr4wAnHma6wABTl38OhCVFRmjTnmZwAOZ1zaYn
zVm3Hyy/mJ2jd+DRKFvFM9BGBcUXYD1E/8iKGw1kpwllhQ0PZoIBAbK+0nGErL7HfAsoFS4FjnWh
+OjdMO56hAoxYjR01yFeER1LMUUSJOs63CbbXkiNWZpKXFmzmUra4WXKE9oB/1lZe5mOKos62NQV
ON7ipMznATd0qDHIUeHSMKmhiqTBf/+HPHro1GTHhHAY/IfhYwmVgDB0OIEDF4zFTHpam7y6YBrP
4msOTX6k/tj6u4Ixl2f84LUTGwpSzlZJgnfpJ27BP3HAlEatt14dFmAX9vAwrfgSh0SfiEOSdCGy
eR1bqLYn13v+RL2qDRXQk8Fdp1CDuNSTnEyrJfn2y2g289TxUD0Erzqj6bZwhMMvhu3M3fAB2yGx
FTcKNBdkJ1XQbhZ2B/ew0tNntAFPZ2E0JZc/0rcjNHoqmeBK1pswB8cLnMKDmWLqLeGfRGIqVA58
H08mue/yq8g8E3mFH5AncZx7ILJT4EAxzO8chmwACVla+AiUeKSyT/ljMVwrygFhPLKOO55JoVFB
dkKigBf0M3uftlYGE+NwV07QNE+R37jAtsC1dYgLnBsR8JgGpZy7U8gmSq2PNdlaG+5NlX9SiO73
qxIMdHo9VBCIA/otEp+0gRYT1IjnAngVfD8TySuewdnONKGMZOdKiJGPLHUQT1WpEkl3SYZ9C96N
5oOwV7wl+udSrdPGa0L/1uAm1AobSFKd479v2GkzBXtjjcataKeAg6HlClIt8Yibfh/lMO2ldtye
lPZRNAghO4rf6e5j4WKrZdOXTG3yOFaOVsFkMpVKL1mVvo/+fEJgCfuHCYNkoy49kzhsE35uM3Nv
QYalup1v8DvXEnEsIOljqf117uuUlVnIPLWP9mpRj57/a98TxxG5V195W5TsuFUS4PZeaTRhQ3qx
kmhiT8HGN3rjYj/o6hzzvoDgXDpCb3yCL+b5wx662unfIINwrkQ7hobagrVuSUbSZyd1eGzZW5JQ
69p683n6dn4PtuUAJlSI63oFUTZY238EzSWrmwpZaNYFlTcGy56yxtiU4b1PYEaAK27t1SCoM8zF
2/19bZWRM7hLnSEL+Q2V2hsMGSrIug7XUuTvExL394i/NYzhdMchk6pjeaE+10ZJ0iBCe7lWYGTP
19aT52/K3tB9qOKuCYiPBBo1i5Vu59weJZQ9OKHwZAyTIdD99jqZyA99AvhUurUFYz9+H6yADruK
SEoP8OEkgYpIsJhWLaoqHc77Jh30EosCQm1HZs7Gqm97H1w8fTj/Vj/YaBQg8zoIo7Aw2O7UpNLW
1B34qKLR9D4+hprXaIGWS8iDjghKbEErq421uWu4Y5mY4g/Hc061zNOOsZadDKosqoMeJt9oy5pg
vVSUym2UNepbOL3WAPzFn+iufD3bF1LCFEeVLrFFJTRXIJLv2nvbP3NyU+8CzUyg3Vbqp1nlWmVI
nX/MyTHvDCTmZXpMGu4M8rsk3p6nyWgv+l9OJV/Q01cF3XY4Y3Zv1toEsy6ALIRv66ocX7RY015Y
G3w2gESyxT8mzaiNbfLcKjHPs2g0ZoxhRtimwYfj2RjVea59ijI7x/uw6Isl55nmRFzJH3lHVRLn
ZlSEgLZSmqlJroYRnZd/7WLQEPghRUuGSGOFEaFMMLfsBwFmLF7vpmpVp0CUlpq5MxG6FDbQXxAi
afkr8TncOnW4LBicDjtoqKYNevPI+s2dxg5xhnciOwPBhayOe6/GGrazqn7TcIauChcQi9QM0IRs
M8vw0v+7Dfo5qbnVIEEqwkcq8QpQI1zDiRdxAs18GWToH0SPEZGWEiygJDFoAwNLjWGqvWh5+fWF
C3rcTWtNGpUn/HzkVNetk0l38s9ZeXwGXU9UEAdSioAlszUflFsoRlDSELtg6A3EbaML+Bbq8uEz
Ur1uT9sTv7Isbel6R3xyAphpJ+MOyrrZQyKGyApF+76zAeNGJc471sLJwrVmzmHmv41Fl45brMfQ
5QasEmv5zi2o461hHZzRQpUm+k0LhNlTfXIolmkZWxSJvvv8HEBw7fDXDcAtYtQlLZXU5vRbOkvE
pdMMrwSFBVIRwfqx1D35EaIg85ohmNqgAa5VmV/VdE8tz7EHAPsmUXhm/+h5iMeE4FEAc+xd9qJ9
qgeFobLfCn1nek8xeul9t6DPdjXvNv+HburQXCYPZ97eE9L8f+P4Zc6FZ+uJd3i1kOutSIlQenBJ
8Nypac58v3dT2B5HDnn2GEovL9l102H5gWAJ6VwIvplT/jLSz/vxbhFmyCb9lV0PVVqn9wV8StuP
5noR+wfU4ocgjTHn8Znded3ms1ZeYY24lkLm97nzPKKHr7EiWVczatUILCgvf4kabxuLPjMypnyT
MMSNeAtvbPLMbq22zMbEApxWyZtwmkezrQuwwGdXanU4sZ6umsa1aulyY7w1AcnXo/msg90MXrPK
x7vA8NT3JFt3ch5WVB+I21jXspUwIpX6Xp//Xk+UqxEIGrq0yV/4SzZLHJ+Wn+HOa+TAhRkM5r6+
HKMRoi+w6xsdyal//0mJlW+eStyOPzzCBdJVGUvH0416cJnMM0VZb7nUvnwJqjzYM8ZFvDQNcuH9
QD0oFVQLv8PAE9jTCDEFo3Tn/EYj1radf7Sc981hopwxv2mDKvD1T2QOG+G2U7T9ourx3SNuzJLq
ftbYof0MfPk29OKQpgkJkDIC1/pdVYfsfm2ZGMyv1DRV9AdGpKtWp/yaObpby1lctX8VDu3swnHE
sgJOhH7ksGOvp3oGKPWUpjBHZoBqU6c/i0U/Noptp0ce26DBVLqVLPC8PClohB28YleQbczbH7nP
yIlYAlfF6rL56AlNzGSrszG3Wj7l2002WKy2+k79SP0zcT6/FTUWS8yRAgC5ocbZmI0cRG1vpKdY
mX6ukl2CFqUaBqENdKyt6sLqj34JP+UOTkFPGkdZZdGBUx7n1NWTrS61RLMv45WeEbEp8zqheAVN
hEGLc3DTQsj/aOPvWdZgbgUrqqTDhhzo3f/P4JeTWnoaNgCBrGqBImeq58lTJH/HTbeakmasd+OE
wPYEDZiVolLwDHQw90KVrhjmelsrXwy2VrSnNWMBnenuazvPUnDYVnvjVjwYAiBfZy4gFd9VuNPm
VsFoMPw0ntAL1JywAxCjpNTCkpUHNNBgWCixfO++i4y5lBqedOoDTNDS/IqPWOSlTszuVEqQGoB2
WoRRdEsYb0qNgUVUdPo62Oobk0MUlq4qcoId2tai1LLWu3Q5lNGvg2AUyCCU/jix59WRe6lVWS3r
kEofVT54LwrRSxYLJtzuelHNWzpjN65/Y/ouyLegIFIgm6OTYPcD7xycIJdsfyW4ROLwjBppSnjf
6B31xNK89UJVhwPcF32dRxnxcRyalIYQFPdjkR8hYLEnRt2sR5Tu/86Q4+gwRnOXVXxyl6/6cyVK
YgcNiZ9HxVmLeQRFJVbaDJW+EOUjYGnBLpUWWfPsuWPvsah9tkcnf7pTBw/qNFiFKc6CyMRLlK3o
R7pPBXJ1wf0D7O1LGXEdAiqEZ0KQxKRiLrejUAphMPwLLqqMnYWU/4+GnMArT/ZMHsv8La8YjO8/
gt7v0cqCyzO0PyGytKw5SKySJsFAxIH3JVdNbm5fjJEKGwvpfH+gj60+VvZPvnMnIVrRH6eM7xyi
TKMTeFg2IVpkktMhNHU92vkErpY9YRdniZhwyFwUl/xDGOUB7WwcLzr/IS0j+7NE8T9RXGHJbGQd
KlRyq4qSn44zmpgs0zj6GRFMu1Of+SCMRO3w2UDHP4aHLUrHO9k5lGsU5GLlHwWg1GOd/VAD62we
zu9rTRJXFl+0rbGdE7nbGyLMkdA3DgS9SG5/X6K2ED5wwfGmlXvdJ7qMxeHqMslwsMisb1SRZFan
aRoSxCVfHb7QsxbfI4jTq4bZ1JqfqeQfS1hQbZJaXdOOnWnzEHqw6oT2gZlPZyXmnlxSdLzhviZK
gcmsbTSSxrq5csXqCFcrr1kCDMqWUb0WZULLAdie4/+yKBZamIohhaWtJdYUGoVrrix87eRavSfG
ufd0Tq7S7+K7pZrw054aOKE354fyFLJ5yZnyIAAa4qTVGW3+ckg/V3XeVeP+scXsdItz0FmLAZQC
snawRVGrbpkl7+n12YmMQWsv+dLs8QeUD/4SD5VMCv7fwKUOVdMBLkpV+OSQid9GEbuSV4cb2D8/
YFehp7b37NSMiAspF9TFL7J1D//52wWkBfqtj1YZNALyHbiUBKU=
`protect end_protected
