��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&om.�'\�Ӓ�G@ʠř.>z�=�/Z�����$J<6���zG�:3������H���]���M=�z2��PM��t�C-a�7|�2�Hy(5)MQ�~t�DBy���IMN�+���ё�&P�N��~zR�Te3-x�'�x�c���T�uBܮ$�z�%h2�X�=�$�o�Y��n���� �@��>��ZW!���-���BƳT�-����:�袼���~'��p8,��+`]�)g�qS���<4}�jԝV�h�C�[ b�����`%iGQF?/��!�r5�)PJ�zD�瓶�yRȀ�^��FVO_�|8QJo7���%�f�Z�r�A�����0:v/��g��O����A�c�x�%5,�KFػ.���a���6�G�a	N�G9<��?�̲d���NQq#k����=��vV��ݨa������\�����?�u�&��G����f�|�i�(�Հ��f�Xˉ��V~��Ø8pwm���@�,Y�)����%%/��-p�Q�`]Gw�f���5-�]U�`6���TH���0}�GON�e�}�=�=��ؠ�N�AӤP������\���ؿ����'�>�^7u6���0~�"}�Ni;Ę���Kq?�M�So�?P�ԴP�k��_8�RH�#3M�������"��i������@mT�`�8>���z�<�oM�gY��Ώ�{Jqf���N�7�{ٓ��,(@n�v��*�ȓ��/�S��]��+^o:��N}Sn$���[�+�����*��d:(��Y�����<e�T��@��3ؤ��r��S^5�$��p��I�?��~��n� �٠�&�wm��Bh.@ւ6�e0.�Ta**YrҗP&g��Y ���o��\���(;��*�-D��v�o������ڪrj"�t ��g�P'R�S�C�݀�X=���|H#7� �$WY[n�",�+ x��)��lz���ޱ�����	Q>��(|/�� ����z�-"��>�f���E���4]AKF
h��#|��5�~���D�'��F��F�4�l��>�!��|
��Ȉ�2@{� �_��=�D��T&b�琴u�E��}z<;Nl��r�St9��s��GJ&��Iy����y�ߤ�RJ{]���E�6µ�N����=���0��"%�=cM������8Ƹ���GZ�Ơb2�����MI!Z�dU�0�&�u$XW�>�*\����!�����-����!,?g"�9`_�9��P�ޫ0/�y!�� ��VtG��d��1,�����
`y޹Ӫ�
V\�9%];��q�������`�� ��U�>['bh��o��WGuFʢ2x4����GZP.Ƭ-���}|=��`D��>=��槔R��-`R�@�[fΎ�aA�X�-�u&ƍpS���ץ|���QP�X�;�⏵6�:�^3_�콘�.�Ѫ����zk#Ѻ�E�EĪ�k<�F�#{��^��Q��j�� ׸1/uqV�<�f�0������;��I� ���n��nŘ���I�1�ٻ�#c0�=j��vi��;x�&r��"1M��v�C�����:��%`	��D���vD�����ѶqT�{�_]��!��cÐ�/�����f��V��xC�
zE��6Da,�E�.�	�c5	���㿤�0^�����KF�.2��������(��T�C��n���I��ۥ�u2���}v�(�v���=��}��\��rR��pN=3�Z$!���L�;~J|I�u\�JP�m	~��'��D,v-L���tk/`r^�S&8���Ӯo�j�8L����	�Al��~�\�=��rh�}�B+3Eg��Y^3 jQ��i�aaB#+�K�I���c��uI"�x5��Йx�!ۅ�]�B�!�0��׭����T���K�ȆO!���Mܙ|p�f�r��69u�o�'��lzA@����[��䆢Y �Z�V��".�m�e���il��k��E�P�hHI33JD�R�Y�G��*��d����s%ŭ!å�;`�_�b.KGVQ.���k&?a%�$���ݖM�7C\.z}���9�+ ��>�Z
-�c��V����aD8��O%�ٙ�℩-�S��Teg�D��I��ޚݲ߸E=����6���e�`w��/o��E���t#���n�8W+B��Ţ���)awA���=�pw�kĥ��&���Ř�A����1§��| �g�>��U"#� 񅅜����/�����$�������?����Y���{��Q���BtLWKӣ�R��t��@�i8[J>��֣�����R�RH�k�ϸOy�\k����G7��}���n4�>�9�'�Q�jJ�R�GI3YmĎ���ý}�:~��!Z^\�zb1Ok��?�NF�����7��:��*�]�,��V��ۥV�j�3�2o��j�;g���C~7-$V3IW�	bS
�#�3qM����g�
I�95��q<��82w&�#�h��\E��{s+���4]Е��!������	������ʊ�Wܣ-��+��L7M�:��J�Į7+����j�S��CX����J���v����ɤI<�Z��r�����ğ`(�4��s��tf^Į<'o�Cn�&r��Ȧ����X����f�:�B����@�|�$x|uZ�B�b-j/���MQ��y�%�p*�pNt��H�*W����>n��5��X���ǻ3���A��Ef8����&/ (������V�����q�l2��5�A!���Q5�	Y[-����-b���8�ܬK����P�"�1�; ��էQ%�0��b�����Nt���V��|�kb��7.2WWʍ�䗧����	��#��b9�u�����88 [���M](�V}|}*�[[Q���Fŝ�cAx,B?麃���;��a�	9>������	�����~�+�=�՘�FٚU��	DSc���
���ފ��|Q ��M>�_�yd�����Y���8�C[G��Tp�{=\O���\�j���9,!2#�ˁ|�a ��s����^��$d1w��ٶ�O�M0���e�"&|"�}�A5��%���n�B�1�lSK؏M�����x����{��D��}���޿1Y+�X=����V�P�o�O��nt7ݙ
r�i�.}C�`rl�l�`�/�+Ҳ�آ
�]�����a����$5��m�p���=��IgL�0WD���N�`[<&"�U���*I`���[�u�a0��W�z(y��W�0Y����A�d;X�i@���h���K�e�Z�ʮH��5cK$+H%/M����k���⩨0�uthԅ����z!