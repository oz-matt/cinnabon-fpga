��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&om.�'\�ӒiA�<�Ad� ��Oo?�s�N���0�@��Z3
��OY�+�S������`�T��M��Ey:�S��#}���
L1!��r]��m��
�8��+(�����d�$�4���ɥ���M��B�^,4����*}[�ȉ[%��Zڎ��lʮd���P !��>YI�8q����A��6h�;�`}f7�<
d!I�UgP�<�L7�#�9��e�>p�v�U��3 X���7�y��;�m����r��<-d��H�i�~oI�bb*ր���1�C���V@+Q�:��%*.���q�2��l�Uޙ���������w�5H�����L�};h��k�6�H�7��!)�7�
_�S�U�;�<�9+��j�ͳt�ǻL���:g/ʱEؗ��(4K����|O�&qy�D��і�i�B;�jfSD�o��V����m>GF�'�w���~��;�v�m1-����7��ŋ�)��k�8��6���3j5�o�(�dH�O���Mv<�|+�p�(FH��r,��IJ�ϯ��-q"h?�����>�@?���&ah%�u�;h쬡 ��g�V��c0�Ow�������E�E���ӆ��Gs���3h���[�1 �	������WW70ʁXf��F�o.5?ig��Q1�]5������q��L�c�^h���)܈��`�+���l>�ʈ���b.�e���(,���_H��MGՖ�ԢV?
y�Į��@	�,D��v�=�=*]���T�)% .=��2�$ 
(�W�a����ke��ґ�;~(�{�wA݃N5��Q�����ʨ���q���<�O#t)Cİ*�c������F��o����&ݤ��;��}���U�b�^�N��P�d����o�/E�P��ʺ���Ma���k����4 �3�M��Ԑ�G�-�k���E]L�(�/�H��]��oӥ�krC۰kmn	�}}��#��+{���]������#I��L4�O�Д2��Qf�1���Z���mra����_�͡�>��:��eDf�p�z[�"B������=E��{��`�
��=�'��� �Yɽ�S��CP�۞�N���z�j��*�ƢR�AMd�1z/@�8 F�K� i<�=���B�����ĕ����ja}�6�Z}�/�(q`�7�Ē�]Uz�+�����9��5��S�<h����H��D��]l[���RCHs�7�\8�	~��2s��KRU��7%q�n� 씦���J���H̓��b��#*��b="����_�܂4��n�-?��S&�5�!����>�*����>#�S��A�W��Ë��Ή�Q��q<��B���w9�g�#*�X��&�6�3ХWh,�c�n�5��U���djf:�f������j�x�-������!�<�«���Rm��+�ȷ}Y�a!���`����J�a`G�V���,A@+����CX�f���n7���gMǕm�v�����
^Y�A^D�~x,7�����&�����7��Ffu�]���}{����p��9��I�:����e8D������޷>��]�xF}{��쯔WBbχ���3�wάq�3���ڛ���	]��q�8�8�p�66b���:����r@��%*踘��Ljw���ك0�d8� �������t7�"g[=�5p��{��%K�_1};K��$BD�O��L^��P����,��ޞb���	3/WJ�@�2<���Un�	�Z�k����� P��!Uy�����"�k/�8�2o ��y}
P����G	��~����]�^-��w߅ Y�^�ne�z��;^��� �����Q�ttI�����|4 ��&�}���H�jsB��0X_��ӆ��D�dC�3s`6=�p�!߃#����\��~e���:�`��=���B�鸜��}�{+ʐHi��5�Р���<��Q��x��d�=-Z�G!�X�r<�.5�R�]!�45�U
��k�fxm���?�b�K��|h��sJ}�p�d����OM�Ā�0�Jqxj��P؃�f�ٟ� �kv�
@[<��2�AT�Ρ�C����;EZ�a}T��&��/���8Ln��%��=�Bʗw&~��Y�ov�1��@��,�J����[
ȍq��c�_����eT�~ ,��'�Y��N�D��{X��c��)G�_��x6�bg�+�"��R��w�"a��.p�g��	=oO��\�Mg��4B���cE8k.?g���x�/<��XU
��,QۜKL1����#��`ȋQHT��3����x)�iIN�a,�����׭y�@γZ�V��s~l�Iu�>&�=5�S1���VLS\���H���b7��l*4A�I��,`H2k��M���ԥ����NV��L�D��>���YN��`���c���f�F�Uf��P�����\V��#�ڙ7�3v�b�"��M��h���C`��{F�BA���1#Vuh�m����D�C�z����P��3�báe�? �H��/r�ضo1&��%*�X7�<�׋ ��c�d�ɵ��ز��z�)!��ﬅ��9��c5�3��{�t	����^�m������>8Y+��j6?���wk[�i8�K��01��e����ۇw��u�u���/��_	�d`��u�N��p|��Y���Rc�} �=͡o|��/Z�arh�n�	���%�h!��;�w�70sFd"�[��:��}-�g�����x��%?��M�E�GG�l.8���d�㽔G�7)�0���f����⵸�$��mU<��l� ���SIE����j��5Х�Q[73g���n4 %!?y�-b�	~�|d�}my
�p���I�&>�MƮ��>�o�;�������
��U�����(<�ԅ�Nu"S~���i���[ə얡��K|گ(&Í.r&*^S�;�7q�5���?�B�����Ѝ���^b�S�?aي�zmY5B�p�&�ڀF4'SSt
w�|=x]=��F\��ø��Bյ�^���*��=�s����p��V*�u�	�P.,��[Hdeqa�zBH�^w�{�cPK�����r��~�P�$Ա�1ze�Xk1r�v���e��~*7�����c��Vك� Y�����K�5@p��Z�RK�=��z���SX�3�^"s��o䳩��5���-y`�S^϶����9m�������x���V�{?���	9b�9k�����z��턮>�w'��͍�k9�A��M��ڒ����,�.�oӌ��$֋��� ��V��v�?��Ԁ௿���V��f��o	z��� 3F�vE��00O+-�ʋy�f�_��\�ޚGq�G�"]�� ,<�lM�h�vFwd� ��=c��`%��&`_Ql�t��V�^����*��k�wM`	� ��1�XZң��u�~{���g*�^��Ŷ���P�I
�ц����������K�>^t�������2��S�ug�s�\qh��_hȾP����G�O�9�x��9%,gCh>����Ҵ���)�f���"J�j���-��k����}
�n���"Ug�,I��AXn6|�v�!�r�h(a�M�?�DQ�dz-`_���܈X�Dy<��cN�I%��&Kq�E���\��F(��RA�jx{�;��y�Y�4��o}Fv�ܲ�ץ�Wl��s���~�C�5���D��1z!7���PNNK�ZMk4/�~�����r�˿�	�LfӉ��ICnJ�x 871%s��3r@����m������$s�ц���>D�a�u}۪��*����Gy�� �ڟ��c�<�z�7}�E�|�3T����:�7RҩI!�����!���<[��%+�������\�"�6c��nCaڒ�,yҔ��'��.L���ԝR��7�~�P��K~[jQO_E��GC@0 �e�c\�ʅ�j:� C�Yl@f�nͷ _��#��L:l�I�>)���G�G�L��B��Y=a�z��a��ǈvT++#�_�0S����l����5anS�y���,���NXX߱y�cR�gX�k-�±�S�A��0�Y~뜳�h!쎱����R?�^	[��T��?-VY�H�C�x�|�&[���8�����
ܑo)&N�B7c����$u�z�d���2����L\݁�G�*|ܹв-�����F��;[��(���8��#uNV�Q�j�Q~؏ڶ���\M��?�6r3c+�y�PwU�A����g,na�$�0��Y�����갠���i&آu�l7 -Y�O�*xl}�J/�'N6*Gz�&R���ps7I>�9�)a�0�7�68Q/��s"�����)&�����8�X
�#P\d�,�B0%�nj���{���}�Jb�p��~sS��b�����z�EֿQ�����8ل��D����oC3��@�n��Z��=�p�q�Jy����qX���F23�	t�_+��uԽ7��<9\ ����n'�8��Õ-=���m��V��Q�K��Q�چ1�˫!� ,/0��GL�7�%���3�hV]ݛl=���ɝ���D��5��~��k���{�=�Ж���(n̸���o�3k\�W���1~YD^��@L��A�4V���m�z-�VDg��MZ�O���׽���� �st(����HOؙp!�(g��D/zݟ@���e��'���)��h�
.|xes3=�q~@�~q�ތ������<�v�ʗrX�&@N��A�v���m��v�0WNJ;M����� �sK�E_/�{��곣C�K�ax��Zi��aH}�x����2.��#�]x��'��7Ҷ�_ ���{���,��,��W�d&ܖFm���?j-�ܫ�_VaP��Z�Z�[L�ˇ7�� �s�C|p%�{�'���,��R"���X0Z��E=�s�#�_DC����.H����+�z.�hZ����Fq}^.����ʶ�R��-���u	3�����;N������Xc�jA H��2m�숦�9��fF��	�"���R��F}ǒ���e��'�*��'�9�9-���x�����綇"�e��+����@��r=��[��f��6?%i�����P���[_|�hj]��a�_3N������`(^�����n���]�OhY��$���H]yZ�"ܨ�c�$m�������A���<���1�|v�����?�F&E�9cٻ_ӨO�:�f�g�:ɆS�sʗ