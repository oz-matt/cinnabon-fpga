��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o%S2��-ÝV�S��;Z�L�|�Q�dC�Q0 �"�a�!����J��Jig��ƺ�>�t�N�D,yES��Hkm�I�5Л��gO���<"GnNJ*�c;Ҿ�T�*�D�(}HA͈��`xa�y�of��)
r�]fE�o�I�'�)�%h���m���j������8���M���V�1�L�����*��{�l�N�6�1<�;��f�=���k��<iz����W�MX1���6�sH ����I��v���h��~�*ĸي�i1]vU'����<ʌ���HK�\�\�a�?b��_Ь�̬��O�#�3�k���Ĥ��u����H��G!�/�G��bn��8Z��M'tS��S�m|e��a5lO#�%p���V����b�v�k����).�v��a!��d�x�����;�%�A�[�Uj�t�#�<-S|��� �+�,�o��E֪����� ?N�&>�	�7�z��T^J-��� x�6X�9��'f� NS4܋���b���B"d,��;X��3�߹�M���C�^�ۭ��Ĝ�	�|A��mU�s��,�F�)$G���~��u 0���H�<'�o�������
�y�k��-�R� �➖d]g�ui)&��s��ֳ�����d3&��`���a�����ҿ��]�v�NM�J��=�iO#X��Y�$�Ά����
�I+n����F����kkrF�8�� -׳����t9��G Ҡ��3�6��o��&��r�i�=�)6~�=��OM�r�>�M��#��\�V�l��//=Kq뎪l2O�۾\�'q�{�Llh���؋�Ʒ8��	����4��4IDM(�Lyw粩�5���ݬ�鷠��L�7����	�L�lXm<e��&��=�c�p
� 1�Yl^��5�ZA����IL�&%�>�R�P9$2K���L��tx�t:����=eB\��^8����Hbzo�������yIe����>�ф��Ej��*"��@���ƿEj��iͅ��@�t☿c���yI@��Z��x"�TnQׄog��W2�;H�(�!!eC\��"TAX��w���z��;�h�Ǡ��r	���֖G�,�XQ�"��:(����a��;��Xgg��Qp�2P�!�I^j>�)�t��t� �YĜ(�֒��&�/0�*�A�!Wtq������>�2lW���-����^�P��j������~�t��[+��D=�V�ok3�q�Q/P�����]�ދbb;��B����[*��"�/�.t������>�?�Yhj�6�7�u�tJ���v���lx��b;�ѓ�����DD� ���l\���k�!��%l���W�75p������+�#��ti7�K}��2F`$ʆ��'\{}���LkMИ�Α��$e�l|y;~:�QI�c�:gy&g�00'�/"���~������m�82�|@O�r�Dt ���9�ݲiNCc_���%q֣1fL�̑#�#t���V稁���#O�������x׬SŮl���hy�J�ǲ�������J��qk�s�×!���K"0<�����B�fZ���+&憈���J::�w7�
 ���%�|P6��u�.�qgr���>+ro���E�Yֽ��M�QY:�����-{��f.��-�?�[:�F[��>����P0�Ѱ&����D�Қ<�K�W`��.�v��ꐄ���K�`���\ҷ}�����<>��d��g�e�/��=�8�S��DFy��t��ǣqeb??d����MU��A�׵��2��O�hG��6@���d�E&��*����D��u���Uꣿ&�=��ҪK��ǜ����ȄI�R���\AQ����j(Vo.-��1���^/{�Ԁ� �s(�/�y�n��<�����0�~�!1��4�� =�7�U�V�
�xS�F����Y���N�.���d�M�O�����SqC�}��"�x�����eV��~TɱI�F���d#c�1�_=�K��aR�j��$����_~>�[/��.5��V�E�Ք%�ͷfD�ץ��\�-}�g�$x�G����LL�����p�~>�Թ Լ���cI��S�N�C��:���wxs8S�!���w�k���ZH�.��6$�J�Ǐ��P�h�2�*�S���\��+z�#P\�4��2��
!9���u�����FΓJ�=O�b�]5ٴ���w ��Bdt��{[h*W|9SJ��t ^���v��/��{��73���i���� �E(�k�Ɲ�:(U�*Gk��O�@()ŊJ2��S����2�`�����%�q�t�e�6�<�a��]у1Gg
�U��Aam:�`�A/��کM�>g�y�<J�;Z��<%U0���� �e���"O���.��k(�=k�� Q�vl�1�3s�7�v}G�u��a.��/���>�$Z�v)����;:B����3U�����1A�T�>+P�]d({.�j�ިV%�j��d�1�-��m����L9ydKZ�ȉ�z��w�#K�2r��������pG�L��Z	�0�`Pu懤����\lNn��ؐ*eM5μ+��*skQt���uxHC�kXI�w���4Ε�7j�0RA¨e�� u�8�K$�[���a���J��fH���E�
o3�/��~�	u$�f��j@],��u��[#�Ƈ\\=��X���G[ș��a�?D�B5*&'Ŧ&6��w��c��ܚI�Yޒ�I� �m%�����ܸ�:��n���fiE���@�Q���k� ·�]Y"�[˛q=�"��jh�?6w�����G"2^�B���'M��.#4���g���֗�|�m�\���'/��Gnu"'ε�6�љv&�X��6�r�kP�܈-o�Vo�	�/K������L�<#�����@��Nm}�?��yo=�2�Qd���tQj�X	��"RԽ��g2��d�
g�g�g���v	咧���I/�d�e*a�zV6�߈#���S�b�.�s�:�Otm�[MV���>������Y���9Y�(^��s�灦���/`��I�rn���P��7���ˬ����؈�мn�%���Uv" ������_>=a|(%��Ho$x�("P�F��d|Б�6x2CԬ�q]��8�Х:�8����m�/J�y|Oķ��F0K�|H��i~���;�3J��=��}���Hަy�z�Ѳ"q�hORG
��8�,̹�dͱ��C�&�{�|�Iզ�;ȗ��'�D����\P{�yl��\:�-F�+	�X��^��g͘���Ziү��I�e��� ����9��0�hl��݄�۬�Ț���_�N^�kA9}�@
I�Wv~㺖 H���Rl���	ȖP������c #W-n>��}=��NJ˽0}��I���R�ۓ���e�о��-P�:�L��WJ�h�R 7`P�v:ޤ�zC�ڟ$���%�����ׄ���X�?V�L��:N"��y�l�n�eb���I��={�ލ[�]?DH�Y]�sO:�������ذ�x�7U�Hn�4\�&vdb����n�~��:�Ն}�&�W��7f�(p�t?~���Y8�ܵ<��d��]?�AO�bkʨ���^���e!+�zRxχٹ�����͌����HR󩞈����U�	@����Z�Ɯ�A���ҐזQSý��c�������?n9�"�[V��bs��6׉�8ԏh���7͹��npP���)� �٩j�����������[�'յ���/�GFzρb�S[�I�-�;+�1�Na�{0�7�����e!�_EG�!��48�5w�d)B���WAvnv��K�����m9^�v���f�C1��jN�_	i�Hf�l��U�!{�t��o�����mM�~���J%�\��d|¾=L��G��j�n���2�[!��]�$,Ԩ���Y��=X�͞���%�`�v�J�J��Ԅ�`�ݐ3J�c�[�B�f�{��<�h�e��5i�L�_{��U��P�̩���TL��
ꗗ` ���b�1����Μ�r<<ɠh���JG�H��d1Xs�Lb*�H�htФ�P�S4,��M�N�S�S�B�1�(i3��Z��%g��|j� �5 ��v�(ƙe� ���L��E�
>2�&�L��5Ua6ނv��+���_��G.�V�>��W���a<z�hD��LG��P�n1��B��L���J�>)�dJt>�
H�|�S:�6���S���1��p�h����
̲M��p>4����)Ib��R��Q�v�A�9.%<NK~��mW{n�:��h��SA�m�7�;]��A� ~{$M8�aڟ����}���e2���%���E3�mt{��1���O�]GV����&��'k�����Qo��X�&om��;8��n�]#�Ń8{:�r�U�\�D�q)�kQ"[$�>04+͍�oƶ��I�*V��RVu�����S^����3#�w����g�Dh%�/�S8v@H�J��v(�c��$!��#]=��[�*W�h��L� ܨ�x@�3���B+���%��l+z^���/+�"��h�,q�"�-������Z�_�6�t�>s�6���sSf ���g7s �5%v
�+(��fuF~�fm߸1�#�z�̠@6	�}��;�)U�2����I����>J�@i"�Tٿ��ɿ5��癑�,��6���Z��}~����}����#�±X@NC��f|"�;䶫���S*L�T�RLR��x�5!X�?��M���+���kV��o���C�>��Nб+Y�:r���!!iA��տaM�w�: 4��W��.=���0J�MuJ�� CP�r��p�&�F�Rj$'6͉p��yڎk�V�Qfbz�<�,(܁W�f��$�S$`�9
�78��b�O*㮸؇���V�|ܥ�� ��B<�=��J�B�j�A�{1�8+k��Ol�K~#��ʊHG�|0$9��piIޠ:��c�U�Oi�'�wĪ�č ̙XCU��X�pþ<Y��2���Q���B��>�ˣR�A���Py¸�qB1�A��]2��  �.�qK�K����?k*orټ�/<�����vR}�k.3�5t�Z���w��� �P2ǯ�3��:����]�[�"5��S��X���玻��e��b-���J�\�yP{���(�.�(���a��'�ed=�b[��'�^!�_�j��η���������TV~��xC
��15�zt1w(:ȁ����9�;~ͭI�6N^Kdw�g@�X�+8�E���[�b��y#�h�烞�~�1H���AZ������KN,��H��F�J���r�n:w֖���LU���2�?�{����^�z�:oR>�0SU��/~d�pX�,)w$g�{���^�_r��Â� ;�yxz���^J�!�$_�,���}�Q4
n���2��q��l7�j�e�[����س�EЂ����%�-��LR��+�M(��o�����R�&tr���`8N
�~�f;S���[�B�Րܣ�u@��^���kT�$2���f�Db��a��-)���Ӥ�F-r�^��L��K�B0{7��Ӏ��:�%�����e֬�m�E�i�_�	��@tR�s��V�N`WF����%5J��e�B>���D�D�}>���]��0��y���1�����eRl�DV�D�}�J�v�Sw��C��yfx����{q�3����S$6C�F)ws�b$�z����p�'L�c��v�2�*���Fǅ�l��ҡB�h�8����h��v��`���xi�UΘ��8 g���F�^�.�*	���Е��f�}���sb����).�Ra�	l@�
��Z梆�c"Np���G%�I8�)�'���^��[���sR�w�4��J��^��7���ҷ��i^��)Ϣ�����L��>���KET�O#s��O�naR�W��f'jv5��r�W�Q>�yvC���I� f��c8o��2_��˄�[�p@h�Y��Tu)2檭�L�%����nT��`
�;>��{T}<l�ahm�)0�f��dAJa;p�".�o�Vg6UJO�eu�ti$�+����,ܦ�m�_#H;g�?�@�{�OD��(F����Z����9ԛ�.%�L(!��G��J�
%������l���kDjVF��,��2�O}ux���h4J'm
qo|FY���P�H�����D:�@(���r+Z�clm�0�b�NI[~N�h-"]���2�h�6�+�V_�`;_�s&9y����Ts���̉1 ��p��ZWP6	�G$ ��Qyg����� �r�t�� A�J��GC��_�C�D�wm��0��_�u�ˆ�-�/bVL����̍��'5�4b�onU�6xh ���TS$��������+1Ĳ�I$��t����-RF�0�(<{���Gu/�̫fR¢3j�3V�1C^@n���y�R��^��A\�"O:�07��[ן2���/�yr�-�Ӹ�'2�5�a!�1щ�k��9΋���8݀t�ԔHG"�jbش�| 7��	Ŷ��!�	Hzu��%RD7F�!��d�r���^�aКeRm �i}_��������%��T:?��Q�#،eq�Yj����\���0u-�Z����]<�mI��2������hB\����]��[�o]g;�Ǎv�I.�i�yDTx����z��x]�<7����+�3{΄�~�Z�N8�aRS�]z���K?W!�Ξ�U�ȣ�8��	l���0���c�CV򁚫��ŋ��9�x-1�b�����Cui��uO�Ř�l�E��H�M�[����C��@%�_�N�%+��)���?��8�L�jJ�6bߠ��P���Z�ə�ž�2���X�Ò~�J���	�-r����J�C�<@,/f�II�`.ܙF��t���>m�4��=.�`&��!��&l-5n�$� �#���5�����=/w��Ƥt��eD�q����U�`�F�w������Y�=��2e�+�O�*?s�s(�����sW#�,V�B���="�1� �a�F_������"�|�f��l2�W����!T=|d����na8�~�ֿ�o�[�tU�f��t&_����·@��X�����9�?�MC�59V��
<�Ӕ�^L>�ȓÀf�E�Q9*�h(V&@�
%w�eI���+f�O/�����H�6a	4�pMF�_�ۑo�O���h�J���́�JK�*��[�{!Ŗ;��V�����`pW��������a���k$b�9{�I�gW�/��0���ٶ�U:2�UW��%P�䂧�p_�퍆�&7����I�և���N���T�jK�+e�k�cd#sSP*��H#_]7tj
D�7�|�����L�w�(^Gu|P�!�X�;��yÙ�=�%�6y�o��}�}�E6e�7�Ch�c��=�3��&5~�S��݅bg)�;�>�K$����W�D�$�/�Q�t�H���O�L���kd�O����5�7X���k��P6���.ϚL����S�����.T۷u�l���� u}�[-�p�侍VR>X�(���Z��|�Č��$�>r�K<і�Z��;��"$�D�m
	9
��]9�������;���Qi�DQ���7vU���s^�$,[<f#m�X|��?�E�i�\��������-�̌oF��05Fy6��6~�C��^�PO�M���
�kn��o9�_ȟ����My�6�w	-�^\3z�RG[3%�%�GAV�d���~�9~��8����:Z!�b�eۙ��ą��V��o�)��<�F�kbs�7�����=�Eݴ��S��J&�4��%8u�v��:��p�e��?�'H�~�A�;����fVǈ�d/�o���i�\�m�Bu.h��a��=�،��+a��ܽ��U)�����f�8�U�����W���`t���&�`�@�['l��H��
��C��c��+�5-;�$ɤT���<6-�����`�t$i]��	DYAUA^���	���e�lW�OK�L��E]�G2�[�4`u��+ʪ#��b=���i�"�!����3|�t?�C�%Wp`�&��v�ԽRTe��cA��x��+���Y�0oC�!��v���O]��7�x�V�ho���A�(���x{�5QT�����H�CM��dzl�{p�b�MA������&"��Ҙ�v�}\�8�`���N��|qc�s����?VSB�?vߐ�E�K6P��N�x��>�ݙ/�+nT�v3υ������L>Pm5�[��\4Z�}���a,P�;� m�U����{���E6Y۫����>�̹�J�/Ma]/,'qF��E�)�*Ui�k�=�!g�m��Rf�rPv�7��K���J��9������k��c?L[�\�0��=a�����S���=Rb�(G�!������3���n�Н.`N�<�c'2~��9�1�����������}~��_ ��26~��n��]�Z���?)����+��ӓ���{h��#8W�C���B@q�`v	�yz�U�k[���[k6�8B����\�d��w&���0�b�Jt��x��rf��#0A���z��!q��*�i�	�^Ӣ��<��(�	����'j���~c��^�S�F}���X�%����_6a>Me��A�
|���-�,,�X�����T-��.t�8P�)�F��ց_���7�hVn�!����{�˝��8 ��mR/te���,��#�v>����i9	��ә'ӎ�#���B�V��zQ�x��]xm�  ��L���`�Xq��_d'�-�tz�IVS�.��`X.@��ʮ���f09`��\��"NC�w�>%�1�'V�ĳ���Ł��R`0 ��¬�XYO��2T���٨Ui��V�9�N����7�߬~�Z�H��KW����ٛ�z�'FHFp
��Æ�B;�t �ܥ��.J^�15.��%�����c"�T]s�]���]5��-��}���~%�M̩����C'�M4h��S�q�n5Y$1��Z�1�C�-�ZuRy�[/e�����G� �bX���Dէ�&�w�](S_D��^�z�� ����l0d��z��bn��2�c�� tKB�Z�*%i�جa{��[�/m�he����H�4SZf�A�cq���,w/l<��BG@����
W�#l���@�
��$�a6 H�<_r���0�8�][�wh+�B|2̻�'��<�ɒ�֋��=��	�NH�P�|ǹ*�l)�%و��1|���9��X�\�}P�,�"�aoS>���l�WU_1�ayo�-YS9�wiL�� x������� �'�h(��l��ĭ�G3/�󁫿�_���n'�7�_&E��4����4�=W�D��C| q�t���GL`����׳�o�_�Wn�#::�ioc]�F���H���� ���Ľ6&6�Lb�%�ڦ\��:TI��M��v��0h���x/������1��8��r��^N�{�֛
?.�+�""��'�'��:ǙL�������h�)��O ��)}¥xT���@K�W;�V�Nk��&cZFv�����6k��8��5;I��~�w�"���I��^��l80z��k����Bo��2��G�x��4=��3Q8� #-�h����^������Aph��qY�|x�����{+ip��9���S�e�� �c0��<��:�)��3����g�.�u��5w�lڛ��`DZ<l�h��`賐K�.i0��c������+8�������T�P{K��,��v��('z��j�³��euQ�M�㋟�G�����҂e��������i*�c�5�|o�R�B��_��#�+Y�SG�}!�l�	�qYs5�N?���(�����ZN
���UŐ!���̊�,�F? ��-��!1+�!9�������Ni9�E^�5��/��ܳc*�=�)�/��U�����q.���8��&f�	v�ϭ�c��s��鷣��ǖus$_���p�Y�Di�+m�훼fȁ�+Ծ��������)<�t���n]���?�i��E���C�l�o�O�e_g[A�V�����JI5*�	�ͻ\�8C���i$k�����z��7\����'�P^٥H�?<\=�;�ǹ�XC�爹Φ��yL5��f��/�m�T[]�Q�{l�!cKOd;���b����_'9��K�t��������Xy9l�O x����Wf웂H��eU؉��m��͎��-yA)F�98F����y������݂Uӛ�Ͻ�qVJ�69��MA>I`�k&!L��	e�n}�FR�(�Čwӳ�D��nmV� ���һU����J��zh
�/�a
%dNۗ-��9�Cj���:��(ʗj$�fl/��m]j�59���ݬ\���v4�4����)^>�C ��E�[w��.J�{���l��	y�tH�!��^�
BD��!���w�LuM3�+�n����������2��.-5�2��S��J�G�3*c|�����S�5�]j#�_�b�c�B�
:�y��w�$�P�\�O�������<,ZF>��&�u8��D�R�G�[�-i�-�j�c�v
6�a&;HCp��!�pU�/DP�Q� ������k��A�:�
K�����K�f�������gB���	3�.�ۆ�]޸j\+;��R�_k~�ˊ�Y:���r���r ︻�B"�W�9�u�z{N����h(���'�熽�O��{��4�� �^�[HpP�qr���3��t:��sO����L�a�(�R�HO7|���&�n8�-��.�"lqC
p~��Ш���/}72��HU�y������a?���Zɶ`U�m�ƣ�n�>�O6i%2*<�DX��$����!�7��|��A���#�O���܀����9�e�ªm��I��M�7}�1��8Y�86�oǥ�[�GB}S�gB��5���.�a��; []c*x�Q�]�Ҍ��{�'M���?븠Qp�n�hh��R�eћjg�C��{K��i&����3�����%%d��[���]e�)A�n��ܾ�A���6Ubk	)X|$�,�{��Վn�zu�x�nE��|��@�����;��]�9 %f��Ԡ�4 K�ď�_�5���~]���ou(��'���j�-�-��Q��n9�!�a[Ɂ�y!k&�����8M��3\(:�J���~ȱ����_�W�o�Z P��K�'RR����^R�O��(:c��m��ꈤ�_"	�x*�j\���������R%��l�����x�ق{�J7��A�zN�)�o'ic�����-���,����L���6�B�ѝ&gO۷�	��E	W#ñ��Bj'���nY�Ǭ�p�EJ�F���8�O�D�3��R20�h28��˫�{T�Ͼ_�n�ṛ˳EA��Wac�Zr�$���p�z�cG�7p�բ)�a;��v�vUri���b^�mp��!O���e��Lm��>��85���q9/>>X$�Om�h ��	jy-�R�J��"��;�C���e���7���;��qQ����h������
�Da"6�>�x�<���w�U�+�'��|`jr0_$�����bġ@��A�㜄�0�~�zg�KS3Mn�< s�NP�hr�u��+�:�A<E���	�P`�o6Q�%!;�-��y�c��h���>��h(�.�Z�cv� pa�,��4�:���tZ��_�]>\	�,#���%3��ǀn��Ki�Z4���v��뼮��%�stapo(}d؝km�������ژ����c	T:����)G�L)�����A�2D��
�Հ��v��=����BAÿ��M�8ӑՒ������	��ہx3�@�����q�?�OF?t'PK�R�K��u%+ (�]��@���k���W��PDPwX�d��N�x��l�¶��"�`!�5���μ	8�lm��,�Ĭ��|Dg2�����NN��9N��X���"\���^�ָ�����>��O-�q#���|w��f���VN?��H���1c��g�y����Ev.�ƅ��O��>[I(K�o�JO�ewA+�%�a�j����
�}ȇ�S�lԵ<J^�����Bg��GF�I ����%�Zm�X�0�m�oTV�s`���%KgB+l��(n���4|\���|�˅��~E�KAƖ$?�%�����m�h�A&;�!�AP�����$�sMpJbmXfӨy���"�6�=�p�R�A���Yʚ0%h�a��4�F@I�K5��mt����G��A|���zy����~�!�]y�ڹˤݯ�W[���N������/(�lA��;��/�4�A����#�״ȍV]�o㞯��"�k�@��<�ȤgI��tW;�M���' v�^�%r�\_�����kW
����1i �9���������ӹ#7����[�
���
���y�wB����Xx�� e�h+��Tܱ��Ur{_��pO���];��^L�� \�#��M��x���(n!Ù&���c�9�0`Q	ɽ�G���y��뀢��Ih�~YA���o�P��2u�9(��Ou�֋:��k_�UZ�l�&[���艆���xcn��?#�:�n����+��Dzvt���p��t7X\:rqS�8n����f@��)9�����-���\z�h�)���2�y�.��B��(����JK����V=g�o$Ϧ�dcN�w���fe�=���qn�/9���C�M��ѷ�"������YĄ��w	�|��˨\KV׍Rau�V_km��ND��Ү��BnC��Ǔ�U�N:�80y!`�FV��"Ǟfă>&8V��!����z�K"*�����أA�6��B�\�ӿ�B��Ok���W�;�YP��Ӟs����3� ���h-[�x}���tÏ$޺���/��t�]<P2\�A�4��#�B��0$�|���@��Tz��m{�b��8��\�S2zx�܇cc��T����ܻj�x�߷��~���6qω\���a�uM�wX0�W��]f^x���@��u�N�����9��(\�h��ө<�C�RO�xF6���w�R^���a<r	Z�]~���VXT@&�y=5�}��FD��F2u�vM'Yq�R���˫�oǂn�M�^}ȔLlOf�\`���o��K��Y��5*�abfǷ�t�k�i�=��):W�����r�yˑSf��}G;����f��"�7��&��[�5��u.�>vr��`��7�8&DBr��A��T4�ߝZ/�ne�,���b4m����p���� ��%�)�{��@�,gLM�+'�����+�pnr>\�2�>���ܱ�C��x�B-������"?��?}��R�'��	�C�	���X����dxc�����}s�0�L壝�<Yx�~��Y��ȳ���=�������;��݊�&J@@��R��N�5,� �O߉��K b�0̈@����I���nm�\'5e��]�t�P����gI�0�� ���ك+�ǛV�J?� ���;��gy���PA�k����].��X����]��] ��c#�W���/_;N��������6��u"�,_�)��:c`��KK|O*T���*��R�-�ga�W�q��,�d�.�KS�bp����˽	�����z���g��>dHҒz)fyYM*lV�mϓ�����^t�&��S�d��k���-9ҽ�ϜΩ�ͮ��&L���n:�v̰$J=v��T5��,��M{�m_�;�>ኌڭf�%~�g_���ϩ��rX� -��QT�|��%!�Vc����G�7S/02]I�VN��V�oBk:��i��l����s�2�	T	y
@2�ő���&�9 ����ɍ��E����x�}����f���X�Y7�u>��lU2,����ׇ/�%$Bt%%���c̒Ql�����E�2�a�ҋM��L��m4f�}U嚅�$6��?��*�^|�z Y?���崊"p��o��t!XH��5�q�|�.��_0��$���-�dѢ�N�V�y�Tb�
V~�F�+\M�v��%(�<S��Y����(�0>h��e�I5�����P(�T�2u�J�Y��Bd�R�)X+�7�ZbM񅫴{��c3 �vB/	��9����X$�)g��{k��;�j��]��쫣۶V�W��HЧ��O�쉣�.59�����}1V=��� �>m�:	�Z���l�������aa�c�,v��f��D�k�֓/O��#2��r�;�d�~ m��̉�n��	���F���s�
�ά��1Kd�V��j����*-V�'�H��[:��Nz<���ʾʗ����Fn�HH���#s�%��F��0@��{m��aR7Y@���}��Sr/�D3'��$m>@v��k�ebfzk�,���k����jς
�}ܶ|�h��05Ȝ�oT��k��i�fv�;r�ޮ�5ýI0+�YWl�?s�1��L���R�V���Zɛ�bX��^t�ڡ0�Ju`�LcAUq*ͬʼA	�0���&���L�v�5o!𳆥�z����Y*������Cq
6�b.wʬ>yB�?b/f�2L�F^c��r�������r����b� �"����<�R�	z����b/���T�1s&b$/BJ	�W��}^�)�W�S�<	q�5�]�{�{�;�!nJ
i ��qs��^���5�+L������d��!N��+�G�y2L����<��,=D<�̽L���r��D�&�+�%/�[��2�c�t_J"�����2j����'v*E�����xv2܏��������Xp�Ԑ܄[i>zG�,�1�1z��Q[�Z�j6s&��ҞO��v_�N���S��������������X�U�W�Q�:��o�
��g���`!�aꦭ�ξh���n$��^�x�{a�L-�
�u�%.��)�M�*���jCù�fֶH|(���s�3���yϪ߻���(1NHc��A̮�A5~o���Y۬�����F�/M�1$�'�c��܉H�~a�x��g�{��%i%h�����J�9���I���ȿBb���Q�.��*�m]����#U�}�wYݮ�X�TM��{��q�7�X�������*�U
@=��*(�",����J��bޏ,�����x�ڹ%�e7}8h,~~�dy�ﱷ�R�r��r���˝v���L�
�Bvu=h�W��-u�Q�	��c�mqK��H��\�E�,S�$�1-�5Xw��Mr���8]]mXb�{F3�jf�5�p;��bB�.!�>�ր��b�ӝj"��@�n;����]yz|���N�����cT�U��a�.���JWp�	`����&���hM���`�X��G7H>UܠK�>�>��1�-v�F���"M~��S熥WX��uv �`q���]�=��k��:�q>� '����I��$��_��T2��gX�I��r�;%ve�n?H�];�9u}n�z��8-@cu:�����ڐvqs��8��Sˊ"6B�͙?�3�q�@/�>�����~3�IĿ����uN$�͋�xElԲu8f�~�)��J�+��{,H�K��62���En�30��tܥ��қ�C�b�W18����b6r�<���J����-a��b�[e�_��G�O!~Z����L�!�sN7u0��H�|ƣ�b�p.�`YS�nq�����AP�k��L	�+�M����ֈ�|!�l��=x=�B�a�"x1����K�����H�6��,��;����ӆ%M�"��e\���E��:	�E�G,b�"Ql�̆i�@t�V�ȼSX%H��8�S,�y� �����,��v���]N.�� roV�S/����p�.���>\ӼQ�o�����g������5I�%��EP{�4ۋ$��X�١�O �C��C�4�n�1�Np!�3ȿ��N���.�z��=��kf���r��k
�8�T�(�5�޸�а9�Hh8��Q��0HZ���(�m��x��6��E��.��(�q�WQ�)�Ð*�~3w�{����eTG���$\�Ul`��ٻT�м���~ޫH��3�/�C��Y��(*|�P�Sܾ�A=�\�J�Q�X�@I�?�T���$�p�z%�J��5�4B��>X��a�n����!���o�[|J�o��B��
��'�,�)���9����#Z��Lz"-�ط�)B�S *���5��C�*~8H�
��/��G�o)���FBeX<|���,�r�}��De�Ď�u�c����f��a��v�e�jN�'.Ӡ<k�>�*�f}���� ��%ov.ƈ�]�|�"�~�d�9ӂ�*�ݺ�`���x� �6T�!>��C��#d,TҫJ [�[{�7�z�z�:ߴ���7�z	��
���w^f��)���+>��o�\���M{��r�q |�7%�
��B������1�����b+%]6Q�%��\��1Эf�*����2G�G��2:)`�����V�	$��8�ג� �40p�\�,/��@����Ȕv�5+'��L�P��T��m�~�u����-�!�[n_aYcE�C�T�9���v:�;Ȇ����0��H�vZ6,��Kϵb�긇���P�Q5jB[-�A"2�y���G����x������E�=��䉾�H�,1%�x��^\F)&Q��F����'�H�:�Mu��l�?(�n��{((�G[W�������j�#�{z�����@TF
�ɟD�e45.hSK�\�2_.����J�$:��������YXZ>v��1�����S'yRA�&���+[^�k �{����lG?�>+)�T��[XX8$lVЙ�'pGc�O2�͜�͖�Yg�=����-kJ�FfT��/��^db�G�8q��|�&����rӢ@9D�yG4xͲ�D�\��m�k�N�r��wZ��hH��~/�G2�[��k�0q5�/j{����,cSUl��J����e5W;Բ�i}�sJ����M�HP0���ku�}��qr��T`�Zq�	��NAq�_��CZT,D�� x�J"lz ,�G�n�f���H���u�$g�W����hg��m�8z91[Czg��/��2�@��${i$e��3u�S"C�C��nZvp[�/�`�������������e��9-�Ă 3�ve�r�J�r��`��a���GX�	1�X�����?s�� p+GB3�sC����-�����JMpe"����٭386|�"�5����Y֩�����cY��4����rKg7$����[�"�x�9��C�4�~�-�q�
���[��)U�w��`<a��?��@�`δ�vÌ����Xr�\X=��`�����y�?��K���ᰳ�v���>�BT �/VRj��B�_B�	��|��4�w��4��_�WtX:�3��t��t��Cd��qo�4��-�'���]����1n/�>����pHBkI�h�Ψ?ނ����=ZW��9�;Wp�����YUuYy�����8]�@��:K�����o�(��K�3��@b�}�H�8c����rDg�T����+돧j�_ݹm�,���$��,ue@ly;s��*�f/����:Xsꇉ"#5X�~GA D)~���f�߅b.��l��e��̒}������k���7/�J���3A�؂��	�4�$���NoQ�����d7�~�6���i�RpN=�B��Q9#l�C#֏��������������=R'!��+����*y�ER���Ƅ�L%�{�$�7����aj�荍B���l�e�)6�}�o5��xP E��~.����<׮�rPv�,+��6�jڅ!����vBJ��������J-敓UM��z�5�oIDɿ{mi�?'*��%!�z�����7�����sC��	�F�M��1+��c������$�:�f3E���s��;��ct���鮡B.X&ڱ��ot����p2d�<G 3��}GfI�b�������9ފyYI���/��_���?����1���
JP)BjE�r�W5��^���Gg�N�
�������{��Sr.;M&-�3��f�"�ƤPF���2Y#b���sTE�Ag�}��'gR8�ꤦX~��D����^����b'��@y7`�XP���]�����T;��+gRyzҨ�C�k��ؖ�6�p?�~�D%c�I�X��.#��0f+]E|�0��Z ��Cl�ޅ����8�	D7���ro��Wh	a|ux�D*���m)��Re��m#�\ ��B°�|k���/`)闑`e�{<LC��/�}���)�*A�����'�f��m�W2��'L��6:ef:�m��ce�����Z(��%Zִ�v/%�����e8�w2+~�.�Y5�(0�lk8�CE@b�+���0�g�������<�Է��)|׍m��;�F�z�»� a�Q:#!;:��ab��d[���{�'�,o��~���0��Ӭ���:�q����^9~E�����}�&}>�Yqq��N���o���k�4�~�?Aq�g�me��D@b���KЇ}<&��ƪ�0����xre4�i��E�]��P`�S,����O����MaT�sZ�'ypNO�=��R,0��f�{���d(�	�X�{���$9�
�6Pr�-�F�e���Y��"�a�_�~Q�_����$ͯ2!5�v��J�b-��?��y������o����5WjvE�0���3 ��*8��>�ʸOhGW'f�"ZZ�L"?X���x�,�����\n/�5Z�V�{��n�\N��D)��$w8�F�fbt�Sس�tMl��H���u�?�z�ݱ�7m�qC!O��oN);Չ=�7^�P�4�婲JWg&8�T�6�!;=\E�MU7ѕ[�*����P��u*d�O�����>^٠4b��$��gaB�'p4��h8��j�'����7�s���Q�k>���e��+}�m��F�r��i��k�<�3�q�鷄�L��)�6g�`ru������aR��NtzZ�?��M���w>ɣ�-ZY+'(m����WHz��AI!���;8���/C�Frnx�59#wx�)*���9K��E�U*c�����|�v�����ݰ�b�m����WL�U7Y �����+&�|C�Y\�h�cv�a������lN7C��b�#�i��ߛnñw�#wv�i�k��Y���`7h�GB'%�>ᤰn�V�U
!+q�vԺV(�{�@�H\�}���;��2�f��M�N��n�!���湪3�[����� "��w^�d�''�C����D��E01���F�(��=X��GUk�?X#�E��Ѓ�3�jg�k�H����0E0�$:���;�u�Ƹ��Ym$ AY$��n�o�м{X̾j|�H룞͛�=�)���0������T'�f<��̛�q:,�)�=�v4u�T�0 4�Q3O�0�i�����(���4�N)����nw/�w�3ĉ����G���?i�+U9���K�y�q�"�G���Rc	?�/<i�$��d*��t�����^��:�	��.nq�i<�,��8���_�M������������JSԓ�2�~����eh�V���D���:hMύ�Sw	��6A��:��2d(��f[b9y�1�1�U=��و,�#O��֘�ը`�\���i��T��W��o$�"�\�8%�(��5:@8^n�FL�r��,�h���2g�o�hҮ_�$�(;�To'o�6��ⷰ32�$QE��M��Q�W��M%�>^��'�����:���.�1iԂp�ۀg��=B��Wp!���ALҽr�_��Lf����B���@M��5�h֮7�.�r~�F}�5��o:H�l��&fAvk�����F2����p4���G����BR�e�����$?i�fV�5�T|��5سwb�f���V����*m	����нOElа>������+�`B)��hW�N�W6�������W馵'�q��6�h-L�Έ�[�C\�����N�I{'Ѧ[�e����M3�+3W�޺�_b�T:�q��G'oW<�[j\ݨ����-���UU�k	�P��
��(,��r��sK��VO�d�@cD�T�bK�ϱ��9�"����ͮ��ՋJw)����ru��_R��&7�QcB��_��:���aQ�t�3tZ�)�,ś��4J�eweM2v�k�v�[T�$��}ʨ��6}N!Zu�d�՚�	V��k��f)献S*�>�}�7P��8y6�%.G~@�oOv�;�*.�x�*���Zο����ڶ%{{k����i����|�st��8\�ҩ�����{�ܣ�8?�||��P�#����Ka�:1���tΜ7��]��\0nI��w�����^E�iC��P_he9M�ƃm��d�a�~�2�:;��ϒzD��D�9�n5�9Y�V��@`�M_y�M3�ې;�l1XrW��-�!:@q��h�6u�'x���UM>)��:%)	��)�1m�x��֎���xM..�`��X�!8(�����1�e�K�Ii*�T�����y�\��M?GBi8ok��g�`-��&������=4,аT�n.ok��H$1}po�Ѵ5'��b����>�e����R�Q���8 ��)���C�o?�;��7��<��Tx���"yt-C�7�w==� �dsm] ��P�}��ě��آ\��(�;�w:%�]���uMw/����)V�BjK6��_�F��dó�Z��1V0�I�]�.�������<΄�ށ�lI��p"�c�t�����p�J�N�w��p��F���_ّo(���Gi�z�*U{ǆ6�-��;4�N��gr��_X�X���� E%	�Yw��6 ��k�A?�����w�A��0�&[xH��8Ѽ|�y[��JZ>V��Q"�{ҍ�@��
j}�{�7�Rf!l�h'�{�c�Ή#U�6�>Jf6�:l_��<j��	Pv��Z�����û|���>����io�Ѝ�SI��,n8���kCj�M������`S����8�ۢ�0�}ؤ�F��h��F��u^���c���C 1�BM@�벎h�"��ܣ��h�'�����Y*�Rν�z��ƅE��!�ZX
�p>p�z4y��-[�� ~�Ѫ��O������Ho��-_�*�G)�18�[��]0���/IHCX��<]��H!2�����pPk+�W+%��L=�nvR�V�Ź����T��ʤ�Ų��GB�ȉF�L�D���Ww��G6+L<��ǪJ����ų%h����KdikH�"W�� I���X�`>1)2�����i�t�p��ߐ��wx��i���WP���/�����{�˚��X�43��W�K1<N�^�Ǳ���1HsV����SD�J�0!���^m�f����8�ͧ/��qH�v��UE�(�C~���X����:ƙ>�!+�^���.|���@1#`P�U�o�g�?Z<��|˹Y/�.�y��f9�"ָy2�����l��}�1*>\�*h	-2�_Ī��O�ny��Cg�0)�Ԟ��F�)0�yO�mx����M�
5@��@=�^h~�M��pa]$F+��UT�hr���2�ﻟЫ�"��K�����T��ʝ�f��;H�DR�E� ��*>�WҰN���[�i8{�RY.:���u� ���-#$�X|TLK
�
�;��	��ɒ�t�ď�G=ڮ����;�BD{kUC�Gt[�<{�
H��d�7��Ț�����-�d#VZ�B{�Ɔ��yqr�o�d�׷z����"�K�m���$r�IFmĔ�3�I7��M�3�k�T.��� ����h��02R�ҖLz�<AI�4��\��N#�y�l�G���!�6���\�jBP����n'̐�YP�w"�d����fx�͢)���;�0�Rǅ����i��Cg�ΗΩ�`��許��6�� �q!���n/�|y��D�T�/�V�r��t'�WBxJ�&/�p�k�Jk	����v/#�D~	 ���T"�׍;ǀ��Wa��[�M�V -��O�*���

���,��Ѓ�|8�_T�D�D]���|�|-�?4�ؤ�̯��}<:�fp<ya	o�`(��I��dL�!�f��".��� N|A᧭p�V��H�����9a���&���	p9<$��D�A�m.c����P]���X���p�����v;��&&��\t}��{�J}��y����E��wփ/<��#����������w���f��m�v��Y���4��<o��d6��V�e�nUv�;̗A2���+۬��t9�M-����@���$Ai�~��hT���ϘY�;������9�0�SCh�FV�>�T��Fܭ��h��(s�z���)����$µ���Z\���-�=�C�3/ف.���|�]��PNp��|U�#T� ��]ܵ-��� �u`��u���}�a���ɱ����V�("nf��6H*v���eh
��n��R���:5�h�0w Cp�D����m�?x�v2t�=K�;b��٬����Pj�d�Dl��j��
~�]g<+�Y��t(���޺��S�&�'�	�mS��qlL��H�}��'Jik�!������9<Jw��0��t�G���Kt!,�?��ƣlSt�OG7��}N��aO�N��H ��"ŕ}���Y�j��ua��+o
�\����ò��N�p �-eCg������a��M=�3�
+9���߹oL�&����?����"8�Ǻ K���d��8V<+¹�8�7�l$j`N���Cj���-���*�6B#hRCЙ{.��Il��3�w�W����וW��q������2�V�#�����\�:��<�M+��E�Rf�Fe��Ts;�!&
��4�S�!έ}üNq5��1#ȇR����Y��,]��¶��Z���.m�\�&f��'b��B��eWfG/N8��]�!�ƭ_�d"^o#o�}���N��ma<��"+�2��;�Ka���z��D���-��>.Ha�\'����6� ��:$�͐zn�qI���Q��"��.X����ժ�����
@[���lH��+�7$��C#��pP %�t�3!R�}����6k�S�lrs��8�����kƴ8�z�=��(��mBH�w2�EY��$���諌Q6;��aj3�t���8�T>{0��`&�58��o����u!kV��f�b���ҝY/���
툇�k[�
���{ۏ�P�n�����
Y�Z�c�T�߅h�$Ӟ��&�+�[��_I� ����ϣ7_o~#w�9��A�.���g.5'�j��o>Y����i���.�z��d8�����
�9�^s�!&(�2�[��sj#9m%�7	����`
{�M����&pD�,��z�g�J�K:u�P�X����Y�>7H�����_��s>¥�W��ﾐݨ�sׂ�5�!��o�d��P �pŹ��@���%��<h�-3�%Lc����'�.^ؐ�]��%��mo������5f�V���?e�B�;3ZA�9�>�5P"2���P_)�c�9�P�=gQ)�ĮJ����������A��m�*��aG��8X'����̱�� 	��u��X3c�I� )jy#Wf��+�}��W_$炶�+��A[����=��Y�lnA�Tr���2x�sK+I4�Ԯt׀��u޴�LbS�v1z��F_�����f�Í��������É��ΦO��g�aJ���)�k�+,�0kL�>���4�:�ka� �)�c�I��Fd<|��S�~��8�Y�zq��46���>��
���WSl$�*M"Ѓ��#�����qD��&�[�5t��ޡD2��$M�:F^V���%	�Nh��+j�1�L�/��ۅ>�'����<S'���o�#�E+˙�Q������j�)�(��P�9`�F�x#��^��>5�uQ����}]��޾v!x�z���-o�}�Oƻ�}tp�C_OԞ0|��o�\N��	���i�t�S�`[�S`�ћ�3���@���:ݐ�6|ĭJV��wX׻N���
�J"	wO;�l��{G4��S��a|�/�'�E[_��\��'|��OJ��6exQIB�s�@������@�9�|�Kp��ד�=��tv����lČù�߫�4���RfU��r��H�V
����+�2���,�	�e�Jʯ�#�?T"���0 E�'�[��́{�NC�  �8\�0$X쭌!� GNM���D��Y�h��V&u�t$�<�4; ^h�{�d��i7��HS��M�� |�811C�@Wt�ֺ/6z�)c���B@�ޢ�ooV(�<L^�1� �b B�h9>���F&�,�-P���/V>��6�N@y���2����� Br�ݿ+:����o��' 5�����&��]�f�,��:Dؑ`�Mx�zP�e���8'נ�[H��t�r�:�A���O*�`����L^9�n���	\����@ٌ0\>�K	G�x]��}/;l�����㰠O�d�wEkxW`i����CH{#���e���='U�����B֯��U?D$Ğ���D���owO��f; -q$�0ڠd��n�%��$�uC������R���Y9!!�%z<
E1���b�Y����t���Q�#	���(~�� �P�pY!��$�����n*�?���MeoC��M@ֹ�r���H���8߮Ѹ��W\�JF�D�?Ir넛D��E~�Ϳ㺟�����ո:#�j}�,t�E�"֭g��K8�ǅ���>}6�y,IQ6ur&#e?���r��eOW�2����T��1/r|�S���$a���҃l�%6�����,vCƿB�h�����@N� l�u��m!I����Px$�k܂��6v,�w#g.��;l��u�F���W���t��a��fh%ԣ jR1���?)�`�/��>�p� ��W����vT�z�MB�a��)�I@<%�'KC��ir�)`y]��HF�V��@Yf:2�]xh-�&�z�܁�m��S�/l�3x�����l�b;6�Q*��/�)��g`�D�6O��` ���eb��9uIea�T)��������l�v��E��'�*5B���i�t�ֽ��Բx��2�jfM5��\^Z�G��Ŕ���VV��pvR
��:���4�2̯XK��������O��1�6�j���v��`��]��E���x����q��%:���s����fW F(��T��:	2?�e_�D�(��CX%H�@�x����~���ݮ�­��$�yu�ZJ�kE~b��z4���z��bHR��y3���}�k�VK�Ӝ{׮��D�nrW���I�<H�Ε ��E��E�,�Zل�o6(:R7=�݇����E��J
�4M��ʟ`��I FQ���?�ߵ���遡·S?�[Ȧ�}�s�cA?��/:�P��o�Z]V3AY,���?��ս�(�<�ڳ�S��f[q+���2�h��ޕ��U�B��"�Hy�_�/���w��_ȡfQ���U�f���w5f3�=�.8���nZ�
�xw�&�g��@䂓�@����LA�|����/��B�S�95���(��Ep����75k��k��⳽f͐,v����x�ip(dr�p�)�tZX��G1F�X��r�vV >H�wջ�l���bx���A�w.3�Wp��q%�g��Ҽ�d4Z��L��QHuƽk
_ڇd��F��,�!?�BF�֩�N�����:����x�@�����u��/o�	xC���ɛ�U�m]hi���u�"Py�1/}��@��~���f��*���Ps�J���Z"L^��Y�Ybڊ���}�׌�W�+�I0�ۑ�"��_�u��b�1����2����������)r�`���"*���:46ݴ�A��{���[c���$!�c�2���B��!��Z}BmM�cJy�E�ho>6����>�����S��	�S[�g\�˟*^����0�>��ơ#β�^�ư���vz欝����޶T9����B7�7��5�h	�v�i������� �t,�� ��g���v5��v\_���� 1 �G����vP��v��u[m�Q{�C�Y�����4�}��p�@Wf�z�nH�I��ʹ2�p)��m�:��Ĭ ���Y]��̵���+�w���?��=��䜫
%[��F�*�r�{0������@� i�\�1Y����&�[��[�V&�Xv��x�<�JCg4�j
�#�&�Nn�MU*�V��n�M*�w;��r�xZ*�t~|B�.���� ̶��\X<y�ċ��v�&��H�^a�؊�ő�l���[�ʸ<��_eËw��4��G;+��C��H���T ���N_&�:=$#*A�S�	(�9�|QK���^��#4�Z���LF �k]!�Y��u�]��y3ו�����/gqA�1~Y�2� ���;�.���OҠ��$��>���+ä@��V����q�?�ފo<�C�np;�p�	��x�e<���֥�BX%v��{�������vw�[+P�5�֤�j��SU�꒣�ʈ2dC���T0�$�Ŭ��@;ԄĦ�'�����5