-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
o2eHpTf/kxXeXG8npT526Kcvkf/IY5Eb+2PLg+0PScVQSu14lh06Qlr6RDjtQkkVAIwuYdA4YzDE
84mO292yPv+PGiSSJZoVeP/wjKvJaRCrtJFw5sgVKlO414TViYRfbsUJRnuqRIKwSCYgr3OQ/1r6
z1yOcYFQRvQA0Vz4hPP+rzgV9ujT2nPMstJApBlbHLDvsNeX5OZPfitA7UxwYHMAy/nZTy3v1qSi
bcg8H8WjkNgOzyv7RCmlP1A8YrKOXZzs1YIM7ZcVmoHzsblKef7M32HOCArvZ/fCj4h2ThZ23fpG
aZsLkeMz1kEnuVg0CAlxfFeIE4j/ADBWK/kuTA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 23248)
`protect data_block
mU/tuxi0L4dg0oSU92f+qQSiGuoXu2ohVoC3C39k/2AcfJgFvbY6pgxu+CoFRpre4eo8jZa3Rjgf
b3rLyGIhcqHYe6Tf7WgwKyj3lldwK9hmYaxa6DuWEzk8k6NsLKfOXo37x2R6AA7pVV8HyiBM31Sa
mRPv/VXjymJeCnBtzzfNLrkodDULOorl+12LwSq+qdLYXo7Q6XZsFXRhFYHEDLd4ynRSyVGnUVgC
R9z5nN9X1kLiV1c/XTjiR2q2b7eSOCmDTrjXB7fUGx8YznbIvatvy4nXePWW48KTIJiGAq68KVKw
iMRjMGhBnXALQ0DqOkGP6MeGlMKfTm76UNlIHSkVoq7NxghIMsYsApIqVsah3Q2mieBOxp9e0ops
/7XhGpNZ0OQ7z/HttX50IOSKYDMHQcY8DvHpyyIZM/vmoeK9LPwXF+THYKWXu2nLpi5l+s8pvREd
dQoEr/DYZqI5c7MXTNVm7ZGJRoIqTTZcD8C6gXA8XpsSyxREbQtJtBktS21fNWdGk6aQVApJB/P9
QUDg+IUjoulI5FD83LK1TKaBFFjqCxmcHmyrlHU4eyqOGiP8FtLuVyU+MVQNt83W69euxRvZFMAZ
Ur9Uie8lopinq1k/UckTz0LSiNSWzNzSa1nsJ1Vn+wwEy5N2f0GkLeHV7v2DQJcYkO3UrZjWcLy2
wzP6s8TVyxNzxnW4Tbvq62PM1kIG8wAw/4R+cNKJYpiM+N0zACKvPxqumyAL5WFowlHDv01I28ZY
MpKsEx2EQtahfK0jYLL5y2a5xDoxjOoS+RLi3h3LzTqHM6ivKW3wgNhpdBXUGtvVi26N7iSO9mOU
Hi0tcY8b3fwEmBpqUEctCWyi/lTtKqYv1vne8mXIzgcAY505AT39+ChkfUqAHzUcDuZXOB3QcUga
1HwoN0DuIiiCt9M6kKB/kf8YuEKvZuoQqkxr2ICzGyrzJS0/+i6sOhWDxQi/0tmutilDeH5Wt6/w
IZI5D3Cv5cBKbtnHmer6/dOvzdgjY7tMnGehqd8JIYGNp74JspLpi1me6cAqtxyCPd9f4zOhxJfp
AIBQqCyViM6YMMzFZitq10JmuSJkTZM9W2GDZfG2zboDDVLbupv5prDphe+7SuOh4JKAdxH+WRsn
fDu+6cKuobBfOtpuXfwxfVGFpjOab5Q+iuwEUZyo2wMBRx7A6+KOxLXezvOb+syrEO7mKgmFGdff
Bef7DOpZCixSd/sPTIIqrknHzJwHKlZJHXNGzluSvzFoIO05XMK2gENOpzFgfalqf8n0lX+EIPJR
G9s+QM1zCj0YC3ldKOBQSV2u4IwhTLRykVIx4wjFdVX59kAFk0VKdYZcNNrqKFYuoBXwymqZJOtQ
BhcnFcjm/urfDfa0GiDBla9fJ0jx9BhNAc7Y63MPBDxr7JPp1s992WR4EalvJWShbeJ0j9tCnS0y
YYABWIgKnuNR0zwKy2j33qPUParQrs+ieHdL35fKRPg4uhCkdyeFZCE1uS0lMDadzl7+KHUFufqs
2782f/ZH8JP4tGwJGFowDpUMxWN/koemLi03BUrnPjYRwkvaUjNtWg8p4bgWyP3SCmxThcBeiU/z
OzTWGkAFpXAox5/GwOnogcNTLyvWimAEh6Pl8ilYah3msmZTaeekn6St3rQ9kJaVOvDuEDQKhqKT
NqbnTXT9ekBgiNDpp2EJyjn+83yUlFFAYhuE27OHXLMd1cdlF8q4GOkfeFndo12nRtRK3r124GQT
bDb+mQDs0rqCwbVVAofd3OmC/5KzhBA9Ge7Ch3Pwl0wOHg6bbgbfVyOJ7aZKZa4MX7GVKusFgSah
aemExVEIW+37T95tt/Dbb5FH92TWbVX4mLJrkKvTlItnL6Y5wmAO51dTtMlEnQnQDEn1b0VN0pOH
2vKCxWGIXLHZzQZNuxplB0PH2Paxn2a/IY+1xvZcGGCSeNrmjGXcoP4Ba1khVJ6gATn9RtGc6Po7
3UQHj0JEI3ongeoHkYnNixzZ5J+ktqSQBnnpk96hHld+oAj+cKsHq/AJ48dlzlVUKl50m68PUvem
H9Lm4RWxpGThJPm3tzrOHfdAooO07SJnbyMH5qJpOu2HxUWPRxdlqxUkLhVahErA1DmGD+nD9jVR
VKooQ/ulh6FlDArfYjsm1kDzMNsekci0yhwUrnpTtV8rEqxwYKaE7JmlQ2xN9FnvhOG5QF2mIDQW
Gy4xZnaqP9n+5XzTcpfM9UgPImHL3qhIeI9hYexatlFVVYwi8oCmpUhmyciacVIYZk90XHIUcxsx
wZGr7nEtfKEkYWk3alw345+H19Kw251ccZIFhxWTUCq/5WHcc0SgwiHpgpLsGvb6opixskZGzblW
H+gOjX0iUU56Yjtn0Vz0LsQ66QTtlnnCMfFR8GawKwIP4ktkA7kQ2aAGv6QoVYj+W9T+a+T0GwCJ
C8ouoDJ0HY2KxrytJmhw64YZYlN/z0ddHAIKzIw+ib3fdjZyo6+GrxGHZS1miOXP1P5qyage8Nbc
G1OdxbgIL8yIiWUzOiNw/tjH4/V53Q/gVchlgZjwsGQ+mh5TU7i9bbjGEeb4bL29e60fEP6jK4db
KL0oBl//gjzcg+OhsztEhSxS16qUEfl73qdk/nWIKtmcOPTzHh0E/u4dXKDevaNXhixeBgqVQQYs
2Fc/3fO+5x3CXwIXingevsuP+K4MGZGz5eKyv1XA14tD+pnSwhM+gGZ6P+w3fm5vU6Ay7bxFq+e0
s6WKhH4WdWY7ibXRr2QsKIrSFNqCRo6dpQZzIpDAf2Ho2mQqLo2blGKus6UsTVASVxjxPocG66Kq
TpwtbBWoyNV+ggYdWxtKcb5lTT3nhZMdVfOVlhZgEkrxc7Wel1eVpXGvhz0J680sGRdUMxE1i3gI
+B3jB8YWvPCCtOBPR92F6IiT/6QRv5kQANIjYSYrui0LXW4/GJvCA4gkURMhQQGFgw7COpMeHpKb
uDXJGewVRSMunr4pAruk0zClkRBRqaBqxBqDHr8GRJHcsZPq34afF2CRnPxiPFkq8ER9KfUcdH21
JlPfPA/KpuTkl3GAsz6EyZWDmBvuqyiwG/fgibUJQiNth9YMKb8xuaeKrxogW34hLyXANqpUwWF4
3FtqxG0odeJp+AWr4AZQdtHD4sOHIPu4RolyEISpCd4m+W3BGbRdJNoVxJZ+XxOPk99F7MEpycDz
Z3+lto9pTNkFM6sh6FSj8Vwcjqv6ePxRWti8vjF6gLxFldiFH6avJ3HKho0J4Q9SToKpxNLX4Hdn
J+aIIgMRCuoBX9KQGXsQ5NxnPcGwY9wDrf8eAntx+Dg7Q+ACkKEtMr50go3CNKkMhinQYGstpLHz
GtR0Gx2zkQqiIvYiN57e5T+j+pygfTsXo8hJrZBObQpzKDwU2JRnhr0RkKWL14FeFAu0gK43jCjZ
+Xqf9jSF0FnkrVd6sDArltWxnHkVfB07InX+JEbO2ErxQoqJn+fBA2hwxoUQW8xNfb0j/Y5HnHgs
BhuNgwA6bKE2wsgraJGusRfnbYGFDTiAzcWj4jghVWVFKapO5XpxSgRplKJtgGKlEWKf7voVZ5XH
4/9nfN5PZfxZHmfM/b0LQt6fEMDnxvAGrEqGPLfcviYRiafTZF64q59BieCTGf/UoBOJYqChuXsJ
eEOKZ/WehW/uYu6h/4vUhiXW9gzsGEkq52Cze6GUllhQqg/E15W1M1HNx6qC55qizJ8xA5/ci6rK
F++/GZlnY8nTUnWM5DxYaOSnc+VI8vqYXm+HiWdvWNqHursaUDMWLxVCjjN/p5Qk9JO+ZOryLxnU
Ez6py44cGyFEjTSEEqj4Q93D6r71Jsvrrp/9b8S9OUO66jtHT+Cpf+R7Tqyp1Y3uV8et4uE9DqEa
9M+hHphKlhjzR2kUE+DXdq254mDiSuSu7yDN4dD8A8G2GdXLmqtTNSM0HUXju5NEdAfzzfsPAfUB
UoORdnn0loFV5Fu0Meb8/IYYA/1Xo39TyGaiuwdE6UKPXOMp1IJgjIp92iK9JY8urIqlgLlr0Os4
c33AXWB4ahvpyVkMuL4jf9XULCwR2i76m05NP/mmh0uBiYlBUoFwujHPlW3jLsUwH6TwUbFHUUa8
Hhuo/BlOCev1fagfuvEFGol34Ebim4HVFJnzT/9kp2mYVBgXBxed4HvW8QZ5Hx0G08YrYBK+V7RB
86B1Lfn16G6WU+bRBMlTymS5wjAegHLvfjVaAwPCVFQgqcB15CEmQ03n3KcBnvAZrl2aJR1cp5kW
bNYmLGPK56VlLhQhA2d/uSiZxRx2FogqIC3bcZqKnRLJFCHneaHt2+RJ5cg9pbvQm7e4fmZlVgNh
Y0BAOhEeNhTRmfCN5sLpqR/QGfQcjgVdy5t3rBEvGKRrAdVlSQjpVlxNHUOuw5aiDmcYkzzBW50b
3WnOHRvxjVC1+ZfMjEeraLo/Nq3iOEPla641CAOocuv/Lfy/0YBBZjmzASObI0ItDONnGne1SIqo
X9OUGpy8G4XrHt5UbOxpzyXJjY+4xmrKFgaahGQNZepA/FQ0cd+XHWUX496xcRhpTmp+LCi7UhCL
a0vbs+kdKBnjubdF1oMsgJW6tIl63Bgpc3xuhMkQeJvwMSF8DLBlrDb7KeDDqWMaZeHRQFyRW4Fv
T2exUkt6xlFU1njCQHAK0jIY361sfbss+/2l6CdqmYm0EVIuxtUKXclr7AsndP8FocUcYRzVkQ6G
oFXIK8/NUrV1WPzgOatlRSUjcJRz9j7pBRDDnbuq9/3x2hK6czsBO8lri0eE+iRvL1j0MBNEusL9
Z7pVgCkPZU1ohu2enSsb2PIKTPbtapKM42aAij0thJ+3PVteLW+4aJnSiCZg0IEpmK4tK+MmwTYA
xUSIL3Lzdkoeu/iVOe4YOUQ7TeLA2iQqLD0d6y5DL3t/OmjBLVwMlw8KNUMmQFBX9qwJ+fPJ7Mv4
YWY6oSubBCirxMA9ORX5FEVaQQlXyp2OuruBlgbN0a+cA8Bjn+/QTnYuoK8ZlRhZVjeo9Iz4Bltc
R+f/COQgAvjff2PXfF795vSoDOj9MAQM0I/VK8wGeE6xxnN3lFCZyJi6mXHdFE1HmQ7cWjtrRWHg
KXozHeXD6+btSChlUH+1KcHMLRn9ImCs6ytDIOEzuPKqQ8Wy2QNf5v2CHALxeiQldHx5oEh9KiwF
86j3xp9jFJkjM7uM8E2lKSIV3smA/eT9CWkuepxXJ2mRQ3naQ38cAupvRWNYYFNHkCNSA+G6zltD
hegjWqVl1bnMWqdFOsgL2JeLU9RYAizn4EuIw6ExFbDy6AyFR+lV5jliZj89KrTjHS/VFLPIl0tk
XJlJ2h8QJ8p+P1k/OgkZv/TMVjvXxXaPf2ohw8l1QfmAgskQhSHyR29YiCx3R1YMW6Jy+JBpUr7L
MSevLBqhGN6X2TS7k6GDq0letdmrpylS3LuyMLQ9jtMAXQJ0U+ff74Qhc4ng3ymxe6vwAUycBSSR
HvoTM1gdSRKSqRZuE67CZ7n68Be0yY3N/ESEZkWEg1c8XIEm4os8Fy/ZIPbI6s6nZ2k1uv1YUkEa
HNaJavfjT3xIKIjprdPh0ZwwC5R1QOMl5ClPRr+C9tduXR2WT2T1tmKAFKbV/SxL7vBY2LdKU9/E
DXM4I9yC19v4KnmQHDJxNchFRR1s3txIuyhf31o2zOsCPUjKeWTlNvt1LXW+76ngYRa58cEHfbGM
Epd2ElpOdEnPJEZ7PPWXIQuabdavUYTV+2H+UVKRZIUUaxeR5A2H3XdMmKcazWs4urVPcRGsyhiR
qiH9cb5BEm7dol6XwTVGazeC3xnSHNDbMLrvBC65ghAMjX7Adj4w8ooOvcANLOdIejLk3nWRmrpT
+GdxEiJ6zgu4ENvGkmxblkqvcXY8iJIBctD3FZOanf5JcokQHX6Z8hzf43rOTh72OESCS3TnnUBX
U7JOb8oQg5QQ1qZ3PJo/9XpxXY4mkv+g1Nc89rSlaNUtLyz8MAHZtTW3PSTd4aIWDcNOWRvWCHKg
yZMmTI0dqA+yOa+IIKp28zn4wN5I/BcLw3dOURWMBkiAQ+KyjKP++Uw1ixmlmXzPEu6PPNW4Nc4o
4EOIx5NnYM8OEQe9CQCNzTTs6EmAWd+RtQ8BrX+tK0NbyBBW8OyUHvPdeLylltWRNILflc7puVs2
4JGHhOeZMRb1H5KSOXN9jSKRePuwwNf7lmq/PDbnrn8PYyVWRLRTSryY6SnUf0zf85OFhHWbgAMH
oUp1de+zcOGG26Y9m0kaiRtEeHcX6Q/gDkPlRBkU5OPxRrZlwbp7b8VMVMNvCB/soZvn+vBJK2YM
PDwDjWkrV8qb9mAadQ/YbkkBvd1Ott4W7PGrCDlvaNAOckY9xK9darYqaZI2HsC9bDiEBRaFLjFb
xe7OJ68xJsOOHp4D6HZw/hGtJAZo7Q3aqXSIRJHLnhR4g7jbUc1cEMgJFLX2vUFXqv7oJQlrFpE4
vlLeoJXrgeO3WtusthinVw8UCA5eAd1y7lgKFI3A5shAZOTTmjKdkVg3I9QzDrtMg+t5yWer5zY/
97deeICO5lLnf+DqOOtCyjz342G/t3YuwLsPDsjV0jO2NS6un6afLk9dzzAiogij3eNTn8q8Bn4a
NMDsBHFjJLPKKH44ZNHAxC8G8voh2SkY28OHYxHfDXCCLaG34EflxbeIlx5kTvNGyKPmfjx2j9Gq
NVyodxtlFT88UThoa/3lF21vk45oZoBd4dz2etch14jFqnkkr6QCIr7gLYcDJguu4ztrAHx5Yjol
ntpfr1YxHhArUqtx8p6AYUKHWJFOCTNYFLZ3pUMjdfZktiYSTatYjuxipaYEPERATKPTW8VX+U/t
+897PSZqsb0uV9YgCbOL4tATZE817TkWm5eQ+rNpGTgRV8HMYkwRyU7up7516oJ+1tS/oz8kVqxw
v+bpvAL13cjhXYesslPX2EG+R5zi5TVFCYQVCgVhkCehqCkaJ+q8+rSEkB5W+m5W1BEjQFex92Qw
v+QazB8fxjaoU+/Ue2BJzjA7Lajz46AsQeSCzkxMCXw5ku/wejt9vhIyBQrJw1/NFenibpIvYzaH
LKPYeKDTwH7waS40T47jGyN/XLN+smU+nWk0tpRsz9jvQDbaIjslQhP+wX6OhOqH7poBU2T0AjEu
ncm33e+3JAey6ZsyYzjlA305XVW29VhU1RBrYZNVJL7WAp7GDq1YCqBTWGCrkNhT9FVPQj4sh1ZK
kN9jB5ZyxjvVTqq4Ud2kXwxXE3Pko5KmDOPlVz8ZbjEQu6ZKqhu0u2lWNbHaeHI1isiku/EuULX1
AIAC5gI9m06o/H8zUyrTprbI1lI7ZZDa91GcBseW6TBeqp+f6ElR8HT0TUjo2WGcT0XMLO5PxuYz
3b5riE7KCT71Y/LCV6E2qod07JVeaZVkSQir6xggbIr7tXVmMh0axSpuLmaajRV9M96MpvoqUdRe
uRMretaFoT83/GBcFzYa0ZnQkTuIC5tifdR4FJWhOw8AIRQg5vgKgjaDxGwrMVTBnMC23WtwYHal
o355ghO40doX3wXNxUc7e6XuIFmFmptnvhdajnIqQcuDRBdP8/XjZvA3lCJzqKHKg3i7iMuS9zYS
mmGHuHNEgBLrXRZY1P8UXQKvik78NgKUN+H62o8R8kYwtou4ULDgtF+JhDXJzNr4UM/ndaT+vMDh
/Y4oI772a+IoOQfUHdrJtK2QJB2CunGjPGSVwqGRng8wDFthJ61q8zx3R0k2gcv3AXZEA+dA/dBf
AcB+RyusmGkoHmxSrNGDyybaezMO4d9y4S/lef6+aTPBUXFBEN894i6DrOpxZ2CIV2+vpvf7G1pK
ApC3qiUsG/lW+8RTY3K7t1F+7aeZ9K8zwK1SG90KeJdLRFF1JFWalKy16O/4Z7wy23fbP9J/H/fF
5LhdZwZpN+PblNXvUzO10xGhdqkX488cYCbhV7+dDX7i83wIcZBLVkudKQE4dfRJuaCFpeZN7u2q
cMjpBrc7KsTZhd88O7VunNjMZx4b/lQN7ry52LaJF8S/MOPAdbjIICI2lkvZIq+y3g8H0rHX9SS+
jiIOteWOTRVEjmSGlsKY5TbVdtqrUqTcYvsKAusxuUVQKVvhsJqRoob0a28x3McE7rsoc0g1nUnq
eoICaCCuepGcOJBXWmPMKB4w4PXgGA3JFX5IJj251830txDv4+IvQMbIVzvchQQL/dTf5AMQmmX4
XpLwS/U1z2HMYSdaQeXAWj2Yw2Kbs80zl860rIwL3shyd6rFV2v6vAXxM/KE/GYEcMHJ2WV2BCj9
rKAuwFomgaS/axWybPmgxWyuJhYmc/nm54TcpQd8RPVQOwUiVpyp1kuqTTFNKgViJrUcwnHrHWXg
4nuujCT+H9wNmwiTBpXq7YuxwjA9a3ugWDNjjxEt8DzZlbExpd1WmobyG3ddpMBF/mL2ytv1edvV
w7MO6NLrx5tP9M5Z4UDTl+VzJz9AIh6+yVrqiNwY6M5Lfa3/pL4ImFEarrzZTobH1e/yjnxErZ8A
gL/+Jcb5lajQOb9cHIJP6HnbmjRml6bW4TTA3P6ByFDxjaV0qt3dQMK5YkFKENgE6rLRrklHl8ca
mLyHTEyN8SjTJT65wgAKev1oWYj28epvjZLxg1M1b7d4ZuZVrwMWoKUUJQXBufL0FfArc9yhVz6L
T10AzgCxmijkF7EfyRMOVc4+8L8EaL9WzXONv3J79RFhLCTe9XOeG3F+6+k83HMM8vdGg7kJfcJv
N0pl5z6tBeNrh+NygEEGlTJhnWGjRZad2OktP9fG8C2cCHHO4K4kbIjakeAkX33+LBQaVspobPxF
t5xZ63KU3ONrBL+T96ITfW8SHRjqUd8ochbaE2mmZOQkrPatZ/qyzFTU2I5hVA8LpHpAeqFzDqtT
vhs7J3qSTB8K/kff1Cw0r+tFFEUd43MX9xRX7PQ8VAJMkaM0vjlNEIPDnR0k5y+euOdzZhRvPtxT
wJ0ih1QClR4NDkfQ9JJakUlmLD4CFOOCX0UXSCf3Y/IiJCGM5/guD2pa6Z8b2c2k6HXCSyW0ysEP
01RIbuKnVpBj5CwSAmf+bAAdLLBjM883NfpRTxEmmj8BElR7gpL7RyLJBXFBuaLEC1kKV1ybGSpR
1RRynVqVGCx1v/4AgeNBNQ86PWgrbIkyxUPl7HTLG0FwAmsclZqsWV9k0ivAjzCsOioeDL8lEyUB
xn88ouYRF9bgvV4T/4zxLf4BNGgGJ6B1S7cZDfgl2Qy3G6kPKx7/+Hs+TanPxVgPB1z9XN4Z9ovG
nDHE26NpisHEGdtzQQkZ3exEx7u+1lma92SqdihhBYEprg4n8dYIugyan5QVumZ09V9vUxiuaD5g
qBptjO3ry4faqZYD3jkvQ/eMlpnJkLjzhQ1FGPEATKINVcEpDi4wwiRIAkSLq6JfJme2+meuDCV1
ZI8bD/ks6YMGofJCgGB5y0p268lUreL/c+cMyLio8P7yGonWyGBUMVyHvcJ6yj0eAPIZjAFBt5MO
lf+Gjj66FhfYWM/DOSDphPijUtOeFmonmH2gWDflWmaAknRH/80aNhjaHoUUefuF4YBCRfCn5Q8U
S5YBBmXveYXN4McvGlzv67hioZYMaqMWuuPeu31ZSsT5fjUBcPvOXVU1k7msIjqmaOo0HuI0jivr
qIOJyCRKCHWsYhMJOF5Op475Ug24ybYBsWbz8iLZCaMITYh09mmcBmFeEK9ttti/Wftu08AEUrNP
nk1uKyzn11jo7EWFORAAcVFP/9EyxxIbvOIIGOzbWKjFbc2Iywcy2x8zPBTvEbQ3LNEQbv7AW+TO
4gvYGnYybiPJ/yOdBanprMNv+HzR9aXTCTkYTcCdbArKOetfYUZAeNnAiZwjiBgvIOFoQtrcTZEv
QzZ+qxOt5DKWV76F70+M3fAAlX7vzW8Rhk9vn+BuzTa8S35uqUil5WWI14+xORj26bYvAr1K91Cu
fIzbZG3aKof/jbmMOZa9bruiozBedgyYLv0Tvzi93h4ftS0nirxWVeSQ9J1E91hKblCQDR8VYwci
R15E/kTFdlIgcfJopN/HAXADc2Jw18lL7iqkrwDeAJHoLLovdJNS5rqXvKdK15VdAZ6ir5hmUajj
0EILchC8ww6+gZPwfzTd47wsivJ+B30KMibaBo6WcK1RcNxO8fCO5ud0iMcugzpvDa2W60c2kpSH
aLjUYVS62vRZT8PNTaw83K3fQKtO1WDwMMNSyOu2Q9coQLrVxGAU7G2bq1MxPHfdlQnx/vGs7KR/
VnjYmHG9GN7/JR7ktB9UAtonEdfZH1PkhYhULs/b0cCK4ox0bgKj5vmTdwwkmL54rulOtqsPIrJW
G17DEB6E0zqk2pnBLzVykbgOtfD7cRzOzZ1yEfwpvYOV0vCXFdpvJ9r9QiM0XCLGLoMQBcAcwMHt
2IUwhzfqz0GoFmnKJpC6vUMAOik25prddYBGKhjAFLW0S0uydgb3UYNJf4qMIdQD+SnIdOQ9v6gU
0lrCJLPb1fIrYZTo20X0Q1hkOdFf04pER5/QjzDkFFcmW/Rgjle7l2sd6/Bz+Cem3cHr4nhpoyNo
xZd1o1VjK5Ua2xQyl18d9X2IUa9XeWh5vJE9Q7CMyVxUjLL9F9dv10/NBj5z2cEjJzxoTXpAJaMN
m2IPJUIt65cPh8y3aKBYCQUn0xSEtZ4rdsWvCObLbeZrj4ptvCD7lbAIvQG5i/j4ocj27fNM90CL
8p6ob5S2OpP5RYddshOedBsgZLeORcA38vsHoVLbl0HRxoL061PBL9YQBYD3QoijBx1RLjlIwtA/
WRD9A1qWCcR8teKbG+lHJ7pKzltnE0dGkOdw3MjGtS7B5gwQmc6NSwRLh7ajZurPlyK6sY8UuEy3
A3xVQuCpLAOJpiJAEbDDaXVX2F540j5P198YtfZZpn8hVmZ0gy8g2ZypkblAHtfSRJaeYA63OK2L
C+kG4D/nAnvBgFyx5jueH1F+BSBg6RI/f8IPHkL6OoOkVrJjjdRsco/+Ik8u8+zwAv5Wm1u4ZCfe
WW1jXpDWiO2yumAzQm960ad9BaLM9PwgZ5lEicKHpp+I3DQeTX7hQBgEOknwwjBS9fRh4zTpKcgt
xKr+ZF+x02UJ/djzS9XB7TNf40vhAmKpv5U52E15Srfbcg7FGd+1IgLQS2gUVmgqiZOLNJJqsWVF
lKRHtSHQ1wcjLwX4yz9ngXhLQy4jref22diXM3ZVc5SQMl59xwf7Tt6PvBZ1GoyQsMnJfUQjB5Jc
GKEdeM16vkOPy+ilT4p4AjARHkq0mWXp7E+av2NhVv3P/yPQjZd41WdmLmOowa3xSHkTLyzVtCvY
wzvS/C46U4oHOnJVbHbM6oc2myK6NRQEK0OKFjzUcMJpAizhx0+2mANFZa5ydn++bsI9ako8oNYe
33GYOohl/e2W6RamwbruEBpkD3aR5ZOTj2CE1nrgofgHqSy7+qa2022qSDki5fWzseoeF8uVBs9p
28aRQ0zPAe9GwEsjmIQoUjSUbX+VRP8O/DzoMEP+1cBBWpvfSRwCglxfIyypbbCj/2eeSMaQGaHO
Vnvpy/l5PgzFhi+X5rsZaJy5QXIt5zgirGjPn5xW+UOnVuhn4F2/DDBGKxT/tWx38qm3H8ZdFZUp
NYwWjka4yl1eTZkvowf/bEK5/rPlC+rxHzGNJD8ebJTKhkCjYUTHIyz6ChDZ7Pbu0d/uCWhyh7EE
9hltFGlaas+it/NhpcuBTphgq7x/VuNUX5rDLB3K4MjlgMdjBpKmaAeDMf5aS/KWnojm5pIBH4mP
EtvzQ80+oOuqCBj9HXm+JDLLszF5alHMXsctsM/b+1CQCubZDredwBL/ryyWh21Yg965RTU5XSog
3IfL3sb0bmsF3p+4asOffr3BYsn5Ng/O4G6oEabxhUWKkS/wuFEUs3nvNsWChjE17fSGNnIhmmML
InGR93mri4z3Sn6EpMMYyVazO/oRk+vtuTxmtB9oC7WUb5IJ+LbqGL78mAU244dO/+XibaEmaveM
IxcMp9Zbrmf+FytY1VViTAqIH9/RGX1iGJbg3jjgctRLuFJwNH4UEBaEu2xq3wWe8bI6lBvZOyND
Hq5KkiklWhoIeXetnoeaO4eCErh+r126+kmQy90L/nIGAfo6mFt3JxFnRk6XtgyK4rVjuNtlFoUj
18yem4sj6gn67GB308Eb9+LV0IlO51BrVuKqNrmXb0Mo9mTaAWJvDMVDgsMq/SFhzTXcbSpMvcDh
nxAQ4+ROistgWcOMy/5kptTw0BHRnlNzx+NB66seqCVVlrIYqJiTdVHPiRaji0yCMgQUEJRYUsC/
h0xaZICuXcca3/xJOqlP1fGIuaXOnow9UUTG0k38hjWIsCEDJHYHCADKVzSpq9MXNVhwmiyn1JVn
78pq4zYj67T/aGcav2bgAPx5DXmdYs4WH4r29zy51jXUjcxCOz4WxXmZg+Q13rThOuXQH4UfKl+5
1Owe0KjHylTim+OqwsRQ3XFVK7ucpfAG3ntM87uuDxqYmgiRoUnWyjuktBJtkP+Xa53hxSDVK9lK
rd5tam3nAe8w7O2JTjUMRUPf9Yd1TniT11IhOEfIl4CIuWLMuz5I/7FzjDwQxqtzIX5BiPQcz79C
3syxcFWjhBFR7mLr9Z7uESgg/5dOg4fzj79OP5f7tUc45Xc6snej9gGD97/a3YHbCL0VyZpnB2Ht
AK0LvFXAXXvLOMVcCkoRnPfs0xney3JFYmZQ0/JowCMKy/noTDBFXXWGpyqP6JIFE5Sb4AMEkf/a
/FH5i7waFBfRPsO/SLZUa4mg9/czOulGkjSyBt2SvPvh0/1Zti9VffJIsJsCVpfNKNkA9s9kCghZ
WF5SosERQhgXp8THMGZFJwc5dvJFwiD2vAVmgHAvClGzn73vasx+CsLKncrwmQ3bx5JQKNVwzT6V
zxA+R1wh4syXzJwPk60G4HjdmQhYzDmKivPGnkjN0OENd/maSZA72Tna7R334wKwLrfU1TGygtPP
SAkdfJjU5GrOgK/JU9PM3qkCDrYwiQv01NohwvmTs+JV6SqRWxmjXsgkQnBTI9/Ak78SfIShK9q6
yx/4WrK7spl4a0iwx2I3MGZALL8f6POjl+3FvBxHxWGTXdLYb5P603ZkfXuXgKgt3OrIty96vpzr
qHZJ2UySoCWTB9wthg71YChUSgmL/k6VDgHZb5hmw3H9eCO8ouik1uaqqtP6P0odGIrjMaSFBl/S
Jng5CjRxYEcLI4Hc81iTuQ6lPAPsh2nz2USOqCVWE6WspjA5v9yMmRRg+4Yg4ME93QDS5SKt/WhN
jT+atq5Bx1h+YmnNBu3T6+1gaQVv9ltMwvsv+K4BFftZbSOcS3qjPBcLbX1z9SsNXgPyrTDEOnqB
g8YqDrRwbe9miQC+acgzgarPEqtMpmFA0IwSN6oen3GKdfJY7IIV3cEp45uyYsX7pfRLak5fpgiQ
ob786xhXGNHqfoIFkwFGPkj25eDc5W0nBKvV6BDXAmNl6WoQSs8bf0YDAYvuz/BYuVfYVxbRSjg/
W3Y8HOLk8uCxvZY4yz7oaZcqYJhEeb3chRu7mAlFawWIREPtxLi87Q623l3XG7YVKvQ5cImiAPrX
FL1ac9GdZBpt/xOBeinFGzzPbM7bG5JP4I9knsEeI6TZBEJs7ZZJf2zYfHfRhECcfYR46Y7CJK4T
tn6vi7OrQUqlf7nj62O5bj555ogBYb+3rJol0EQNVhH6U5YcGfuHCElkv0fTFyF45Al9o8RdGpYD
nTT62rEHLwc2otSVYJ268807QGrqYbR3f3ZcjFGn6S9fVS4nMmtIm7hQbCCaLWtQiIZp0xyJCB9h
zYf9yy+7xLsbiezhtFJdIBb+s4n9CmpCeRS3hcALKXsmJrgED+awbDb1kkvSQF/TD7SpyKvLoNFX
yd46g9QN+66wJwXEE9SxcuV4+zZ7fQAfioevVdYykySTmqedxUPXxMLUCue/yr0MsVVJlrxHJI9B
gBXyUCvsAe7oyXr71D7XfL0xThujtGNOQe1HRt79C7OCKDh1hqiFSB7IKi1BEoHNe71j4iIzmfq2
d7yALWLozOqMe/7HOqAhPjir9TnKfUXO/4RnjZd0sRa3115fRAazehdfGfofN92kNS7k3HNVTF2X
3/XvacmrEk/OO5X/cvJHn9h2/ciQqbf6XYRLNguF0vilshkzp4/nRJ75oICt5sl5yAGGgkf58Ruv
bsjmtBFvHtvTdsogyGfM4GS9oiDquXoHHV+aMm42mSs/Ux9Dob7ZwuGL0npNYpfWWz6I+QKBn11T
ir9CDJziXSQ3Sfq6hBxE5ZWP8VTCZ+ypYL2wF8E2vyVp/dFXXcnkjEiZlVjfJtGCLiamcm2Zep/f
HZ9wWyvHRARTg2dBLorn/x+xnPwQ0b4iRetcZwV5IB9CZ8Mp7WphwSifdmIUkK85QlH3ojZMgImI
NP0c/xn6CajrAUoJgc2CunMH8x+HT+ei8Xn1egI02XhKaEPQtvdeWcqWlcX8NEmI+C0Eqk9kp6v2
z/zI8/aKJNE7eyOf2MP9nVt9VULkl4HO2V69Qnvn44grHVIl5R8/VpOnLBDyQSqdRKYm6VXFzOH7
MIAze8guJdn0ysJBjvyykF5pJXKj5KRW1NNHittUqDp8EkDHe/u1jtEvL4DoYQJrGKmDXizdf3q1
YGqq1KA/p+vvadMMibZpGXcsIBrtA2dueWq6ve7TFABKWcMAOyHPRLOJYc7I6S0PjarOsbZygZM8
DjobVIr9C3XEytkEkMAHdOn9MrTyhjXqWQ4HBwojwo9TzM9ck0+6IaiL68mejCdgLyVjQ+itgAuD
PBswAhFqWwR0/ja8N+xl5uyYs6dZavUNzS+H65GtpSAzAhcyejWeJXpi4mIprrmlMCNyapN/SeZ7
QToPhP+DT+IooUPDw1qJerWK+qdo69liuSRPFLiUIMpXj31UXtBJ8I/a8luwLPiG7mwMeQ6tguUn
TFYT0zKUzOkYUiJJ7fFCRLQkkFrHrziXzl01uYiP/kdS7Q6bHCbgqUoHODeMt+kRsM22tGoZ3TH+
F8DOlldB3JlAHxHKVGEnl5OOIDQevUdGlIU2+8BfsfyqDwLWKRBh6njZPqP6q1X7l9X0vtE8cNcy
AWCv2Y7gAXGm/wSH5U0/Ne09uvYFdp8PGdX0BG4i4+KEOpuMYpvkZarWmcsvdW6VHLdLr9799V/J
d8AMJje4J+1Zkav4zh4v1iFNIe0qkOowCpw+dhNIfi1/DZKu2zrLdW/cV7nOTwM+w2/yxd832oaT
1kOrD6JYWd2Z+JdzJEOEnHVnGflXWVeTUBuq02mUY5Jnq6YqYqRpH66eQ/jXIIzYCHV+B99hZAU0
t+EnsnXEVMTUwg07A3PDYS2hSYVq4e9SXWkRZM2sQrJafzUOG+kaclZrp5RAmYu6Jm2UweGW3Pu3
i2V0XO16QNBytulYX9kw6J+pwfhtzUNMJWy97zhB9n61nG84/VdMzla/Br4w0zkThDI7m7MzMH/O
NyJPk2T95+iI0pdZW0LPcaA3zPUPazq95JJyqQsO+bQskhPxOU09qHQMe5JvAWFYhjg5wn57ZINu
3hyFn8wwb1ZqelwFsEAej1HazJQd83yjCyQBufto+QR9nTbgpWXSdgbUcbVZ6QSajuUQcilxTzag
XGK6ivb1EWH0o2QnkNFMqLM0KxSRg4gCqqUvEW9IrAKc4hTgcKaZjiT7owZWb6RGmthew2UYB+4/
s1Wb6co44zFxDCtNGp+p4mD9wZBz8/pW8OjHcn9ddT3wiQV6y6cChaOQzBJP6zQJ7oF+G35Eilc4
++Ty45a64jsozKOeIlgaJcHl5/lFedTmplUX0+w7V4iFSA3pqiAqUYrzE6ENBg6sgIqHwQdFPJBw
p0wCz3e+VTBTRiM0krpSfmw3/FVa1F3HgkJiCnXS3tr86eUM6nlKPSGszvHOwrhAZkwdnEvmuyH5
SCQyMBJUlbmPaazrxUzw4cdHusxLAw+yQwzQKbHqrqUNSPbGl5wm0Aog/JBIb9SIEOrhYX+M+FoX
5qdltpGKNNTI9f9Fz7VnCmM4Va5GUHDSfqLP3n3fmyw7Od+r5jmbUY/ACxnx7HW2Zr/j1VGBg6DB
sYHaabWREz8WqRNjEKhEj/x8YFzG9NZTfEs+e3oqHfzo7odgV/rjYe0u+ePuattWMDeKaWptrt7w
LZ703eoaqyvtIZcHenbz3RIXSYwZ+bWqWTHBXH+3d5AYYDSic4pmOx4yHzhc+8fP2rFVEFiBJaub
IJG7BHqSEQ9BQOabACiv2rV1hqFRMyAA78S4Y1HYqSvW1C2pJ7T1/RC6YrYGFCa7yGX3zXmDD2eH
77m+lH6pZmxjcayRonZlfNOFYgM3xCYxTJXAwxWBJPY5ByyztBCiE934L1uaKDwsdVBx4+12SMSH
n8kP6SZhe5djT47zLxLJrOWeTtKgkAXvAKoW8MxZ7Ym7wKObqoYQEg12WLbwIyi3B5WGQqO8PZlo
d3tFXP7oM60AlnbdVgW9eO2L5G0iNJXF5SQ0QDXi9s1SX+pJQt1zbXOYX/QR4UXEyyHH4Ii/G6EG
n7269uR87styilwh5B+n/ci8B3aDhr/WPuHEGEKVLQbcWugrJVvQmebr1V23VGjY9XyFIZvbjA02
lVzH19j0f7tQXBtZy5qd7m/eRRwbkhC63XeBC4I0nOFTMA+0PKRjagrhkZXY/cffyr4LeewxPEpb
MgIaya8pos4HCdJr8tgmFckDpWqOjb7/9/SBe740n/S6K48SMyOl9iTGuKfCDTQTNmh7LUyOGQQR
nX0i8kVFnbAK0GTLpa6UN8EzwiJUEdVb1/HrhEtFDMFO9gFYFeO9jgBLoXfmhUfntxOfss9glf7O
H3mSGSraRrC9+6xmkjdbgGAf55P+sJf/NpkgcNj23sfHhbn/hs9002O60bOfRHUkcw1D+118auNz
eUSmeSOGtE8wdIfK8Glgw5mQLKrKZvtZ1QaYtHYa3j3Oqo/e69b14fcj6JteBVCh5RyUMZB6b+HP
H9X+4SWJSzhGP42QT1JbG06ByXtBAHhEMhVR3Q8c1koWwYgVyn5WT4rsYPX69CJfvqipg62tYmOS
RnfSueQXlLmKZ0odOjqkmwlQq3rBkbjDUg7OzTtCo2tw62ekrylxTTgIRbZ9E560RBjBQX32EkJL
FXV4aBP9DZwdthzKlLYkDk/MsRKEptRMs3mvMVtT4x/BCg0BwrGl4q98vZ4E5FxYOiewaM10S4tJ
tygrj3VejS5EBkOGWe7/XedCwX28DOV5qHFkAmolPB1iHIzJLfxqMrzJjIfUw17RUBfA+SAAeWmf
W02XrnoPVtovnT7DDU1jdK++QiiIUweg705AlYJmQLmCch99y4b7KYFc/4mIXS3GMv8aLy/7/pGF
opZlMmkmjW/dVUNfBPfvD3CQd6mQy0U1cfShX6CHLI+My9Li3m4BNRLbUmsCR0LY7a09+jLSvBIh
3V8ZoRTUYGKwHr95T4KvZVX9xti9/4sMMDLosoasSNh1vdqZzNqcSSAwUgey/DCMZiAkThezdQhf
nLvMcNg1TmkBG307JYpq0SaHt3iIi7VV7al0mebxUgCmKt+WAAIH1QtyUdIsY689hEHtQ3f72/Wo
ZF/bDQLNBzRQJ69N38AyS5XN1HQKTnW29vhdlExrEdi11hBoZv3DGPae5parZynPIczASERLaXrT
b6rN9F/WMmU+4ke2Ge4KCs8nsfyhYURmlUFTSJcfbdCqmD3Ka3aRmq/M1+XHv2T4xa7EOVYtexa+
T8koVY1AYhTT1qeqgTOCnugHbPfRjtTLx9pcglJFmQB/Cc7DU/ENp5EO24f0cluQgxLnNiLL4gcv
BcY3E80tS5n7hkaYT9vMAckQyeZQayZhJFoekYYzJxTxWqS/BvcUEuVTiys9XU1fzpsC1IsQXnKP
2hKXRWgv63Riy3af91HSv1bfvk0+qkFrsnnHWkYMVRt61joy/k1YwYL7dvk28c9A6C4kI4DmmUNO
6wQKGDL862oGpFZAO56Vxv4gEDtY39Lxk7ZzQAJu1/kkL5iSPidzCDSHpOA93j8SwGn36Iy1Sd8V
8DND/kcPGjPD8WUBZSi+CGKrcKh5Uowq4x8ypxc4YGPjl3gemjwFUOA7NmtqKjrexSYjXtPq8Ohs
hGg1Fj8Kuz2x1lCRv5aWXIfi/S3iUBwjLWWgT6tnTGb8XKPUZJOr/6tq5M3h56q1+u2RDDL38rjj
dk3pGWdtkAkOBgjHEEFwA8fHj9GV/MUky4U4WVLb7UzsQInDd7OunEsLiDi37hz8XjKBeHuIW4B1
z1CXyx7cjCPCJa7CxIPZ2gyzMllBCV1MM6erB5YxjR12FszNiimjUARDHV1xLY+NeGnZpJuaPmNi
wv2kuZ+M+7KSRKnIJy+Fzj1tr1v+WlZSLRZ3pXK3vkEpoztg9jctUDTlYmO+B4wCmcRs5k/4aSKd
HKIJIEBqA78louQKzoi+yMFcPECnlnl32sYvHobLPvQSrNIgyJw2ONdPZ6lgRI/hKfgyZI5kP8+Y
J4Er5dEo9UybDMwGIdJH13e6NfJ3TZCzKO6Vt1l4UEkp5hLOUKc1k8X2tfTyz1nZC8Kdao4RAgIR
1sfknwY+c4JsFX8SaMazjsU5UZNL3SydUkG5zNNcVo032T5JTzkdJ8Jo9OiU3uwy0mCxPVadyM01
aiFBWDGnN+ChVd9eoMaewut86+rRQ/KOz4h2c/jaMh4ifaLG6jQ7ohDGBEb78//SezNLQhvd2N1s
IkDcAt6SR2+bPlVUSzeTWvfvev4O1x/cbIxCuLb+5aafSM4SxZ6ZXxT9u2hY6+UpCxNCksgKIoUh
m/SR5FKx/fV1VVJ7MtK6ICqGpxOkcTSZKPNrzEo7FC4KuMHZONJFvR7pNHMAkL5DsvAy3FatHAoo
XWqMnVf/HoQaviR2MLC9Xgmj5a9zksJzttXD9D0I504NICl/AqPDWDOI0mC5N51/CLn8nwZVzd1j
SFBxqyMRix3hnzWIkPkvsJ3Ce4m/8FP9ZBOgZWzFt7yDeDuCmYcAWlfLxzJl3rqMHUEXtl/dUy+w
/SC8EOZbCJxuW4+KvIq5Du6B5mEk51LLIguimvGZRpPGA7IXf+ksYEr13tQoyeKdLSh/oumyC4Qq
JM+pjFKMQ7agr6GRADg9PS9I+d96UQp2JoWt6qgJRbcxs19Da4G18o+cdl90Cu/359VKjff26DyO
bIbtpktWGcPFC64ULQTw98MjIJY0CUXGl0qDJZy78c4jAxdg3kW69wG6R+HD3ynEH11CjUtbMJ2t
nC1ZyTmECNx7IvxnqU6UD/xmDBx4azUC+RT527xhJ1qmguXF7/mP5I7lPwboBMaVGqAYJ4JdeEWA
GxIjIpjOtb9rwOmHRyUPAxu2HHdSlEpy/USGJxdJQR0bUr+buh67IRAVSqfyLUH3JTsuV4frQZUo
Q3SHCspJl8sGZmR1K/7hw+n/oPk6HqPqoK9X3HeCj4F+3UnrV/RTLnQOdthyHo6RKsA1hYUP11Lf
3QMoQcsyQ/wewpyW/7VC6Wk8hNtZuca/f9YugrU2E2AOOF2jqvfw8iz/I0gkLW+/H29PJoX49gfK
6nLA5g246YRfdBQVa1ijImqx0ZN5pmbI2LToWa1k44BZFBk2LXD4/8eKnLs+mDQrYMg0mBtq7Vxe
kZtJJL/whGOofY4i0uoHisMH+5jKkpW7T9RA2oqXQlX/3SmNwcsEKwz9sf/+G9g+KlFqoxtjxjzY
7dA9HOIvR0ehueM7vVABylx+ZFJbaeHZxozptCP1tL+GBygpQderpgoGAKZ9Tmncm1NqUVFOicMc
WgX7dulGnTbzs1jl43lZG0fn4YVJkaQBfm/7O34iNaa3ykDfmkUUDX4qlM8IMjU73Bd0SpljSF6N
8Lc6e/0A2zg/tcmiM3oh3t1btgc8FJY5OuEw221NazVCZkTI0Ue3RgmMM96lVNnh1kvZdILmqZvH
BSnHR6rlMUFC6IGg4rpSKYHOUOhQkylwRuL/Lj7cQ0Y5PbzkZm8Feoeu6ZjfPJa7B8loIJfxAmNO
HDN63Sx2IxUWfXNEpXTlyfyvGa5NE+5Nq3TGxYHNQnzomlMBttP1qx+mEuwH+wQOnN5Y9eGFhRgB
wTBHF+qKvKVzwPjQKOXsZQyq//ww3UMzsYZNDghF3rRp+2koCQpEkAzdgsYMLQnO/5I2VbGWmu+8
2rJi95hbiW1Umcr6g6WXVAiIMlgBjW+jVVdIWxkoXf+pSV5PY93OkmB4OxPOPQg3psl21ueRHp1q
NDBOJM8hd1Cd7fiN8Cuvfmzi8SITf5TgNFnicyOWptCuBbvArY71dHMdqt4F+9Zee6mQTJZ4S3st
FYhl4/CMhhTOSjqtZYePIwj0PCaCijtE8u9bSBspvKhhwTOyQNTBosDUJab5VYEQGhdzOGRoh6qV
KvROwIlGutlCJ9fg1KGhyNWwC+WMu9TsxI0M5Z4Udca011vdLeziY10DBWBFGBkQx4MSW0dPoYB5
QEFLHrcksbdP/6lYquV6rnt5L1jtXf4BPZCwzEfyP6v+0Xio4E9jtJMEmMo+i6B5GQDXuS+TM2LA
y/St9zluWMGxBVkiMaNK7agdZvgXidq1paQrOpV3xhspxbzVpPqQOEZUOWdLi4gweRorYcx5rMD7
cUGGaqbH3S3x0EZBlxv6/AMrA4h1ORtXjGBV+Dp15zwOx4vsqLpmygzo6/rdrr57VKwMVpMYqxxX
yR72rDx/M3dQ2tJsPsDfdXPawhrjPrkNXaHp33MjWF0Gc1/NAVhkKbPUZLH8aWLsHPV/gnsCHcYX
l0OQkE3qM7NCwXvcYBLDtJn+m1q0DlAA3hjFXZR1nGbFux2yB5CqAXZ23N7Lz1bTQjGtgJSSS7Ae
TCxTEiU3NwUU2XnydCY1eSWOwzj6FJUgdP07TrmLH1FunmzAgnfACr8LUm106QiASKw7T6Dpibr2
9STDlqCfVHgz6jYhgaPJw62X3QWdGWgd+jCr1dLxqvjDVbW9D8CRt6mABH5iSH/6b2x0tO7So7X4
HwLJxgvvmdFwwxEb3n+du7K856U/vAKaUNrpTzuhhmQLrIQgvBsOHihHlnr8nZQy1dAQL0Xrath5
mD7rLEce4nCyF2L/QMTIuIKovNvMBbf3O4RdTWhA10uFmixh7yUOVptwoM6b1AXGxyz7ntVI2Khw
wKO6t4FKVyF+PZIC8lZfRYFqA9Osw3LWRogzVvbT1S9MJMjT6oXVh5N8WbxROuW9gv32ioWqNlph
r/tQIcs2IKfpHiSbmwRKVvmN+ZcziH3g3AbtSatLVhzSYquX7WlYeRbzasT2HzNf5sgQ9Jp3gyIF
DgElI6xGGy76vbOwI/q/NgGkllYZAflpsISlrE/3rIV7cdGvgn02Ul6j8IDLOD9EhpAzfN4G+IeM
Wl62k5aZ1r2coCwUutqwbljx9WqGlXzYsZbJrOxur6svtu2gquJ9oEZqjHFYTf3uym1Pq0xv/Mhy
DiZcUbBbadI6gFXI9VHWw4FCYdd2Z8z6J62bfMhEw/hBkF+KqMtd8z7kxIgoANFs1RSl9aFyREkL
tqfjhE87Dece+teYpWzEBiwjty7Rk/lYtIW4bBomt8/vmwlfn4308yV8EVH61FF4VtV4Yjl/n04k
acmjxROg0gPCR7O0foatOzL0NkTRnOYkcABfGCPmNAHZHm8deE8odYKHqOo1Z2+lXEZ9n+i2TZ4C
M+8jfb4FM/USsAwsD64MVbOMsKzPtpSJvCziyDu44QlVjDFc+Wt2L64zpUwo3nUhlIDsXdx218Sb
7RwlxTedQluR8Kmz11oB5Ebg6sRjc/K/CkNaw7/vAQ7xb6Qn3gKLaHtJDdOQIyQLZ54cnPtbNtFa
4sj+K/z/o015xy95aqpFMIMk1iv/1NHzuilzbsPppL6rsAN9b+CMCtOlBzemtZUWGkrhTCZeM5V6
HYeLp4S5d01O+RMRTmz0eJLbcNjJ7e6emqcifkUHhVjlqYbZuI0+SLVYGoTWDduXGSlFm7GAJOWb
vyABZe7VA8emEMJCUGaMB+djsrMkBNZW4gKwrGa9kWHBhlvv20FYMF5JGvwl1aKX1QHQ7dm1fx0c
tPo4T3IvrasPpggojF6Y18oquVsi93VU8Xu5Qy5UsKbS47Gv9ZAM7yFjj4yArkTS7mLbkfKfPXl1
n67g56UhkoWjAQ33W3zslV19Aj5jU8glLGd4hSHjhxBb/dvw0t3ctn8WNMeHp4o8j+rI/ZufQ9pF
mS4Ka9odUkGa3XoBe/lhv48fPonzMoQq65H0RR/3IW9uTjzvzltBu9TLnqrDefwW3krFcI+dcxmz
HkvRLQj5W6TiBxVw8MCCqvkw3TJpJBN4lqgU+H6TcotUNutbkzg6EQc9x7nllCMIClnf5zZTu4Jt
Jgbx2XMzFaZ1zNZrl5oMoAMR8C2HoG1dJlocmakKatdmfldepwK1VlZ4eIivK14v4f8G+wRUEoiJ
1aAj+rTQhPptgPXuZsiZtySdMQRbqsYeigSl7OJYBvcNU28DyqW0phCgLAEdjrf4h8+U8mZOs/Q/
HFWxCEewh23JK8jd404bTkjO2ODHxS23Mwj0q8My3kwRfn7X7V/CP2hEjnlfg8nZXkGVFzvOwRj0
HrpETIBcSHN/EJe7nOah/jU9qlN4LBGdMgpkr1/+Ceu5XwJJNhaHFgnXN1mDYu3BK9AZM0bbeYzN
gafHrLJf21ksEBo/b9bYCnrwbres4oF1YxD0ttKX+W70dUZazUYC809nzTYIi2MTdiYW7Lhrl6v6
N0xmLcaN5HXHi7YWLUZ3hbho+peVAD8H7Qegh2OxvG7Wl1WKVy+QokgBRujiyhlcQj3qS/GanuoE
Hc+RJpA4P1hyWijc9ucTgHvyeEBxts8vX9jjTJZ8hi/zWGqPkWzhFUCej5GRLuytfCe9dQKzmH3i
YqVoZQoF8ARMqZjCxdKgdwq/tOusDqIioPN1znRzsyRtljJHwRyEBCbBcI3mmr48ORLUKTBam5VT
v1+d9XXoEjPdvA6JN+i/5d15z6po06K5GDotJrFXC+bq6YS65KKXxao8Ed23S89dn5Eqj6o+HaKF
T46JtOClIvO8LTvP8CAeRpyZWVz/yO9No9Tz9AZrn6UhcX0mUDiZGVbxA/6BcGTn5mxph+M7LyWE
f8pWFhkPERE9uot+wcRKcFZt+x4i572QbtebqYv/B/Ijhw3258tk8L04j7Hm2/1SIoI8no/6CsHp
FJWqW6uAHCO88oiX/3UqmxR01tTEGny5tEzXf8ehgJVU2TzJObTV3s5YkGboDt9afWdO55rtUF1c
YLZ7og5vp9EsUXaNFpvbTUBQtG/KFbEouPbX6iWhWeoIeBZDbzsawvR+J2/nFelzvkXDziSok/C9
G9C34Qi8IaK4QbHOomnIZkhCvmNHJuCKvHzqKGYTkNUK56nq5cJB0SG2uKm15XjMvgZnhzZIzwJr
rOdZ/3YjnQVCalpn1HqHrNvLKTrHPqHWJoBw2vxquu1tfXEMSPIA6oer0ELnpr/yvNzc8BbGEaGP
+DR+yqAbrENyW4nRclnRewPeCBB0cuR7pWOEaRn34zZnJ+jbbrzA83PCIxFOw5ouuGsmVtSH2AeO
cD4nKhuI0IDiEQA5QEBkzeAe6gYFXFTd2XjWrRgM05+/rlnRMuLNbps7vB0e0jlf5+tGQd4KPnR9
xQMaSPwvyHWZfPZqjDSuGz2Bbzt+64wt7y9eN1zcHkxj8bVSwWK2+VgHr4haB/UHSR78GHo5f8q+
m3j2OktTv3lahD/c8+3wSuRvluMtS3FbpcreRIEv7Wl6iihgWwvDXm7RWBuf0EZ0Hl3xCbbYx/v2
/wOYtlMRSwKHHujSfOR16ccEzGPz5FvjQyoSpCez26pw5EQlJ9BtDh6GoWntKF73JPh6QjpWrVDn
R7nfo0bSIecriJpOIsTWIy89HNvpm/dK+jkKZ9LmdL88zJXfnBkM6Nu4HKGr1gePS+94q1iA+vo3
TlCaEHJd8tE5C1oyaPuZBz3sfxZN3forZtYRsamxLs9uTdpDMhJYS0eyczt8HfPgRnv2ClIi8GDZ
z7/y1su1Dri+oBlc1qXqkIVnddgVJ3i8beO8t8ASm5sRDDc1G27Hm6+4MNADJCV08SuY3ehXTlIs
J4fJdtPZOmDd5ubrf92uV292PlH7U84aUeosGy8e25RZRhhpOG3u+0m6nv0ETrrUMzpYYJceZ4u4
sv114lEXjWCygiHxxi/R4y0wE2OwPUvIIc1J3GHvFMco7DGKeBxxbbt5VjNo35sJaKIQqDNL9gdc
4T1M12B1hIBxaxJp/pNz+7JBMv15KjR55WYWFRz7ptYV6LiVCQdrubucruCU3Y7KkQpBYjGrJ6Cs
0pHVjfcqcIsetbh0/o0EFlEc6A2ROAo+1AXV3c+tVTACLNP4XaHkSTEgvVrQuQOl75QG42Rxczx3
hlqJyErXR7+AkP0he4UgenL8abXKO2ZcqHQ6LCbAY4Eiwftdup8BpjfySRiE9JQWIK7gMcWJIgJA
25/harVyCqUw5PY9asdGccrQ6Z+yKfK0ndRt5+oGgPAt/fiWG+cDcvpEV1Z3qD3Z482tWbiAGDMd
WPnmvAF+JLi9Jqsfaa1Q/8LSTDtmz9j0HOtP+v2N/W4sTVmkUfpYdNhwmeCSNyurWVOPcLxqDOgN
PzLLGdcNsmI++GVkwiDngoVVbioOEkXzTAhDCVec8fojYQYFcIeejW/02LS0373D+EPBw1YUIG/k
FCP6FFNGwt4zV7f/qwOAPdo3mDFd6iXz7nK2QkS0RGrgrMZV+Gm+torQSCAsgIaovLlB3A7D8leY
MdxNEq8G/G5shKNiIz1SMDvThuvDGyeADpm1RTCDJn2BP3Es9lK/sf2ShE4mjRi7B7E2RqU1tn24
L7rSdu7KTHEuNQMP8WObKJq/gmdV3KW34wp/pti5UagEHxylaE+w/Jb7HNZ6TidbaoaJ1H+/Dc+r
U1kcZLqxEt/aqXXyz+nnWb5ulEXE/IIayQrAPWAzHykWv20sGvKGu6O49uQXjIUTk1a2+wK63rK9
OSZoSSLQKQnBHacUK0pHOkc7FpcRHiOAJMOQWNeIWtkXc9VMbOD/JkaJYxwFnpTkROybpCdSctvg
F071nfnUmLROCzQ02qNCVDLJswi31SWSorDbwob61N2r3mxT433Kh1GeBytzwkwxQPNWj3q0q7Do
HDlEwqXwSgNYtiipTGxtlFdNT7LNOAVar3PUF20BO6kkKbw3PTLcKRNw8Q8uWJVxQyup33pRTpD7
z86f5cjXOzvPhKrX/ufahLdUp96f+3gmCJhLWKDgL0OCBWu0lXFkPmw1aKJURyi5+cUUicAeYJ2H
txnGs3lDmpvMO/iC00U71A/0BIsLxXLRaKM36FlBZezOYCWj9S/GapNEWNuWCCKtLIF7+VE7+Foa
FNDXdF1IL0TlBXrbc4lLnSko5fBaFBabs5xV8LCmk//1SCkMDQD+Anh1GFZZqD5X/P48j3nzit2U
PRA/cq4K1v+/FiSHUSH9a/eJCaAD1RL4YSk0ELSlZy1ZoCw5jjzDpBeiL/OERxHppXMACtWOqACg
GzTMHvkYfxEXCgiTv+En7itv8b56YTLTYRHRUAu8GPARXXWkQSmUqRxisLshc/R/3inX36NnfDq4
oNJOTk0bbxVn4I6ZZ90iAgXYZnnMFsMHyqRvkCL4TX+Z4VpL5I4RMQYAp5wLug9p+OhpTi18wtSj
GZna3L3zeQFlD8rf1mCy8x6xGSjyfj4CvDBsNh4YPe+CNJ1ZRelBQjsIkUP8B4ShpuWPTdTstBXw
xn6gyur3v0y6kGcAh3IX4mGjqQ/RtDhXKlejZVa8hdosGRIG6esdiGAuRC6Rk1Jij3JEnDSMf89V
zc+QFdSmZNhsm5UbjH68uhf426NUoIrWQE4Mjer94O4LYZ+X/1Ntyy5mry5wLxO3t5HcXVvH5P1E
wc2IYT91UbpjQOBXpHgOdEMfX580tNd4L6IvdR19P7JjyDBbDED9zBvoSQeAmgK6TJeevo6mH522
qY+cylLd3P5pby0qa9fbjAz4nmcHBxb0QqCvz2XO8syGmQJ8+HsALxEZoWEJOMbJEjWnZQ6CBAcA
sR44iTmDTLFcs5/Vgaokg3jOszPtptVLS//H3V7Tfw4hI4sFOgd594siR2v9yoco+PsDL8bH1hli
7b4h+PfyJe0vNwiIATXViisNWinfqigv2dfJzjpB/Kr1YDIWQfeZhKO3CpPEK2lqf8k9X2ppf5Rk
AMtuM/UzzzfeYpoyB87KSLcRcEGTCsIKhx7xP74Mk8D9xBW2hOk20z5sh1nqsK9QgMa3DIu4BkLU
gAe4ySn1LDjc/TaK9e8EQ9dvXbMQGaE5uQRtWH0kwWHUb2iowyfBmYLpDmfU3yszfWMejsN96zwn
/ANBSC5ycWaHPsqqmlHUkiETeWrvQK/OtFFlodU7uMyea7HCBbZ9jpRuxxUJMELOuzyKQxvN1aqU
sWe8dmQX3GL9TooOXZCz8ZdE4E1avI2PKvjkErOnvKAnX0jOu1L3PrjpVKUPnSH1Z7e4aKqXu2c2
7c3VbDAN5Vp8VwmmSlZI5bMMkFquQMeqrKahLuivvTwjkqaR48FPKw/o5E+gNTpvQx6kByKDtk0z
FzshrWiyTVLA+BlMFha4Zw3FFdrNo+blL8xBUeOeaZH0njmBH1xPEL8oSmHvJFL2zKvx+zV/Rwtz
qgDHA5cfe+JrrUOW4G6iLO2a/PYbG3tbWfKr7UgFx0K+aPeIkR/DWk0uvZhTc/WtYqpRZcuJDdj6
EUeRT5+8WJRjnpzbzrX3tcN1DfuTRR3/9MAswDO7v0JNfy4RbsFVzu4kSVEXc2cUbtasnMnIIhil
twHtln+iMUfXhtHdkpB1Kpf9JFBU3hH1ibVgy1vC8UWsUZcUSZvBgjIsahLbjWEe6dMNnIHp2GTF
ZHXH8kDS1ODZhKircpeE7Sc26uWPrE8yfyaggVMwuKtlTyDlJ8Ck/elJ42Zfv9M1+1K5Usd0UcYL
TmtG9LiuRFHh+uJNOxbFLQYT/wrQJ1wJvPtuv1DUJKWlp25tRzqyX46Ch1Hva4OSS3UOKWhkNXPK
OLXtSZo4uMNrKWS1fCcXh31qW6/satTbYwez5i3bPj1yMoap0hlBnTFkIO0ySumwSjqQfVuJRwAR
nVA0frYEhRFGcTNDR5JrEfv9Lm9owhYb0xCyG3P1nCT2iaa+EaGdawXvr1w7YLmvCt+PfM+EMfTj
hSg4a3aLs+MyoJf+ubAgdAPr7VYVQZ1gMZjKwRwKg0+s9IAYA5doMgBD6Zi7fQvA4voP0bsP9Lxs
9cBjHFf8YFNDv4XzHoo32e/aSRiAL3wi5Kq3TQCbfwjgN4Jnj2iNV1ScNm96uCHtDM4+BZXAPSek
P9/a5kfVHMUzdO5vkBEl9tLLJXR9eW8P8ArKexdJUpwbCJ51GpwW11UaRQsf806PK7WutnZElYox
NAI1rUEKjR3uFhJZf4Qe+byOVFq2TShdjUP4c6ZVFw4mwKFlxJAcr3fnWGaBy3iffec6wFGZto7i
61bHLHKw86i3h/qt9wSwFsD62VLRKYNdMsyZmm3kiRFCfyhLnA4DGV/qxusWv7mw4Ie5tcgiV8H/
ajBWOSCd8BvfjdzQ+GrKsPLKiNag1p3euR2nqnnhGCKWtFLc1zz1kVdSpT0D7sEtFyQXDJeDy1OK
xrgqcFz0rMi+v2ut0kb0ASDQd1G1+qKeRmqrLObHAYzD9gISXZuRK0YslBokue2axgXAqpqHk684
EtPzAT+w/2LH5rZjm0ON4GDHLqFkqsWSTrAVUsVBY+UROuer4JfwtgfSLqd8P+O5LhKxgKukBeZ6
AQVRxmjXi2tGiiFJPfzrtlLAGPAGSJrsiysckfJmVbP/fX3sG0n/O0Yg3RniPUTM0JIY3YIy6DPJ
Ct43eH4IL5NafQ36R9ZDHTZivJz2GGZymD+HAqGMBKYJYob3H34v9My+kQjSyqyb36+FGplVBCqe
5AsbvDLokz8qmpi6N1VJXe73YE4ocKuXlviYoj0pqSpSc6fadUMf0LKHNEOhu5d8XgtcNuZFwe57
0X97SQXRUIkzbMHJYyJ5G/ZE0NPkPTceb3e5DJmv4I3GJidU5bJm/GuY9UPX+KeVDkVYnxxkkA9o
uBkFfKVIwVyIynujTTRkr/0oIopZbqW3zsEqWKI/LZWXBsKkMLeHSfShhb2npPJ27IfjsoTvF7uP
i1XA9daZG/BpsfNotcEgK7/FA0XZ2Elnw+e+x0mQ/yMkdzsWFZyAU3+GntWbrokLnKCXZ3BdjkCX
0COGV6ocbs43zPYSpGk05WQlJi8NQTdyJDs+Cryv9hwl7ldAE+dLeerl5C3D3RIUl+uJmCDse8w/
rMqsVFnyErGm49W7TEW0yIhhQiWUTE0aKQUJVueu6Ma89h2sOzkreIqZ38Zddb8diBW5CIZFNjkw
Gpae2Y8gJ6BHVj3TPQ6CN70gtaxbmWxEK2RLynXRppUXTcGZrjZrYR+iZ4kJSPp5kKjTRQ1kpds2
+Kii4gny7/ET38saXK72Z7w2yDrgCdHfZPikeZiwptrgrMiezrEbhwcDy+ltmyfvsgxkxMg/1GIQ
BCDWguLLJGMEr4Pveke69cJH3Vr1c5K0aiKsvWm2TJWhjiOo9oco/BqSpWc6V5/Fk8C19gJlq2cL
UAWOiu8TtDmsPUVnInmVx1E1d3EYuMuo4UOBra3l6LmE20nbs7N9knf+ywqbz/bciA/gwdy2yO4S
WluQCBjO08A4vabI9Ef6s6gPLvkFKprrmQ5ejA2AyW9nNDejMsNxlFrpJxxLtUo3Upw5zEQXLGwl
pq1gcQXIorxsSfLAXkvEOC/svLErX1oePMQan9HWZcJ/fHlN1Xz5VWOIsVj9ywFEs/4krauHqOcw
TZ1ojY7k+XZOtjk4joom/JI4nDcPaoG/uXfo13FKN1Wz6ZiELUSXB01bsNn5Tj3+laohEuGR0V2+
O7blxnv/FMXHKoeY0oC2YMUKbKTUuUM+H3UhtFubcJRTumP8ExTDFV841fwlJ5uzTHD28c25jLxl
HOkkGD19LeAfXYLnwJzx+Ix1zvAvFAZAIQgW/kK57yTeenI5+0hIBsLM2KwKB/vBeNLUVkG17/Uv
H96MoP4boHCYDv6jr0FIOh+mrplUJeuFz0KJ7SScebwbaExT4jsiXCd9rwI8xgPNaL1ib7qHZSjc
f/44Lbcp7ckDqc01x0mdIx95usgNbBpE6zbmBNd/J14wO/UqgMox1IjJDEP2aiC7Rm8QjlaERYZH
R0+P33EqKvIVG23LqtSLfs5PjkFD+Jo2CuG6Zd8Ty6BhHlA/SajApyMzaYbONwdtMHE5Z3t1REnl
yrHXSQjPTD9rSVrfCsv1t9r8Y1bWbj+6PxjDZUP6wBh9OUdxTfAYLt1IxVJRYA8+wgdX2oJfAazB
uZlVV/sA1RqhA0HjvYi4275yiIX66q/std6jYH/DzBI05iTXsz5/dl6SMtfwX1rancYPZPt4gSF2
v5Rofou/PNuaExVKxlAlqNkJ5s5cAMPSKGWNNu6h8kP3/R0+wn1z8T9Q6erAjo+bb5fKGM+Oq8he
d0dBivxOxM5V0k3ez8eixcB3bfSbCQo/XWwH8BgRCAVurNGUBMiJmISDKjK6XwTwf02swXZSWmqV
TP8tL+yEFODf2d93vHsMa4nyqZPF5h+O5oqx7xW+7r8/B9UhBBVENHT/PxArrJSXAl75riInXsoz
1thgpdN3hrks9avcsZSGM24ixSaZkeR5KVTW7d31BbN0nnTSVd7gvwai4ieVQML0tmnqFMBMep8d
uDtHByYMQvKy7RLlXopnRdOFXimMjfoJMpmD72PoR3S914qtVahoUll7Bt3ncpEO+qIyon7lxNmb
cB+ird956I8UmxrVhnTBXqy8771noXLfAM5IBP15clxrc9TAcGsXj+IAwJ41xm+quIsHOHWnH5aT
5o30YUt61MwUTaMKgallW4RY2weJmrK3WcxbuBzDZMt9Yr5gNGukVzT0pIqqIxRrZ3PY4NVtImwk
MoO8LvX489k0/TWrbB/CkC2vx1uEygENEsp5efMqY6gWqZy+7HIq5mhXHw/nK+Ls5t5IiF9jtFu5
Gntx1sxFnyV5M2vvv0AzzZfALdD6SLizn52REIleOvCG6wmDyer6A7uLy/DuIh4NinjRZtX37mRG
IqgLRqqlYMU/W2tL/FpDsHdURv2V1n6M/nGghI0fz4OGHs7fHVgzxJxBEdMY7pzBJtsL6d81yA4z
HMq/dQ8X8PRj8nAk/4N8JiUfSFMTLC8yGuia/vs685x9fO5jifpJl4z3jLDG/XJBkhrQF/swYnb2
zbfO2DSrA5y2g16OOeYg2Lo+0pHckm6kok2UiaDT1sBeLnOPqwA1OA6wvVIePB9cobCtpqFrenb7
Tfltf8YOAtg6TmnVcu/wlfnOWoC26Wvez85v/v5wfucqU/8z4UNMEQRvFRJuBmK8fUTLK5QUw+hX
mqFdvKS1Eq/TYKMLqEs1P94xW9SO71CwrJIPuLKCN38PBkgJnG4ahVwAJ3cc8NWzIa4Im4BbVxNP
YYiEsUF++xjVgsQz9xAPVhf16sxRn+joCrJC1nIBVFBb+FD7qGRESfKqTJP98oT74xKPip5kfeMj
jPfio0v5Y/Mt/ykfQnBn8deRt8IUKo2vWZz1CJxpAKQsc4+ZuNMbyOG0Qt/Zi9dt7gpIRoQxcL3Y
3ztR3VrE6uuAOCjjYfzR1JWp9o9EwzuNo98/N0+R8UBwaetLtn81bBdh1DVKcU1cN9PkilrsFiM6
8EpEksZuD84NCZIPcXxmjNy+ZxIcJ2MAJaIO2X8XSomRoAh0OGohY4O+6F6nEYGjemhISnw23sc4
+tvd/oTVoDlhwQkh22h3P/cFmxSIHtPToSUQqq4DoiGxehJM2Ajk0cANu8oCy/+8xA==
`protect end_protected
