��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o%S2��-��.���(��D)+ΒP!�tS�~�Cөm*.IF�B�Fc{J��D�<���씪��%7���^�Ʋ���\-f
�*�HQ�M�m��usV�Iլ�B�H�+g��g�{ڜϐ�a�d������D�F��#�����0�X�$�M�Z_P��h=<����<��>\`L�
Ѹs�i�^�>��8fhs�����l�!np��]|A`�Ocߛ�f ��3	���\!��>=$�-yk�M ^h�<�8� ���lsG���,����;�k&K_�����5�r�vgM?(xA�5]V���9	&x����Fi�_�8i��Z�Kf��R��sv�ƶ�cz���I!��$�{:���Y��د���4�wluwv��m>}j�,����_(��gq	���˂X)�,'iv�,=BI�kɃ�E�O�M�+���k�'�/����w����R��(P�V��=�Nqx�2I6v�A�Ͼ�I6�{�����Ү\�EMڭt[G1��H�����ǆ`vpJ4C�}L��+�bN~FOrG;�h��/����ج�D�4K��pR��>'���̩�Q8��*F��, ����1v=J@���}i��+�1c=,4؅��G�bp��Y�<�{�h�6hi�$��M�&��G2Jl��4�/�h �=*g�Ё`�����+�Zjuۧ���ib>�i?1
��zE�J�6ʡ4�P�s�ߎV�ĩ{!H��(���9��7��/��ɠ���-��U��X�둨�y�Uo����K���h؏�K_!�s��M�v(Tt؈y�_e^e���ғc�첁���!�|���h�O���5�v��ܠQ�\p��N�G�i�k/X!��D��tS��c��T�{��%1mmE/}AS�摏��f�\'�a��)�q���fްPM�S�A �zg��\�Y'9�g�o�m���#�8�`����*��?����|C��OXgMR�þ���0���
~Վ�S%F߶r\���W�o�Nw>�P��?�Cs5�Y��9��!���;�>��k�#;'vl.��&�-o�=ܣ6���NFt�Vt�|�<ą�F�r�j^h�0��4�b'����v�=c��d�����5~?q9Q^�jg�y��W����F�z�3	��L&k ��S*ۘbMl�[�wѡsbM������K~1�� �y!�HOP_Jo��ls��6��ɤ��[�v�!�q�����0���&�̕�?5��-w��_�q3�Nx"�p�$��U����r��}�_Ȩf�7_� �$P��!����KA��m����<��Q�-sPi�QJڥ�4������#�Af{E��t�$ 夣�� �GI��08�����C�Y3*��p&���.���S��,}(V%�yWr%�n�|tl�%"}�Z+X�-���+ܔ��K�Ű4����I�9[B������F(�(�nt��141��^f����T��ٿ�izEע�َ��j��M�X�C��7�<��A&Z�$Ձ�^�C
�f}�J�����/46ѵ%1�AW 9���]�J�����4̊�D]x�5_�bs]�.���J#,b�~)�3#����A&|���V��c%=��-w�#��L���j�f`� ty��#���Xkk}��n��:�`C4���ՇW��~���g�U�Vh��*�����3w��z��a��z80���&�&�" u���^���C�׵) B��F�l��f��]�`)8q]�B�S�0�`x���#:	��BN�́�1e�";�b�V�?��r���l=���+���rx�[I]����㑘e#�iw�h.���$څy�d���p����C_��,-[7!{��bG$����5���奔�6�48�q�<�\��DZ:�5����cf%F9	��A�;׶JED?1}m��A�E�2���/�1��&�.��~���5�H$���3�h#�{N����u,$�h����"��+�A�����h��me��vp�Ǽ(My��	_g$��=�-kʧ�D�������(��p�E/9����iv��i�/���:����a@���_���$���N�ꊃ�Y(��e?�T��l�<�4thw��tIx��O�]�:�+���s�G�P��-b`��{��5=j�}�,H��^�D��~K`?���^�*����f?X���a��#��e'^6��Ȋ��wKn}F���A�y-y���*�+A3��6�!|��$ ׼�l��B������9����>����x3C]b� ��p������kd��ܐ6�d��k����͒�ۃp���.]�C�ꆀ��V�=�	�
���Fs�e�@4۰��u��t*��m�{��F�e���V)r��^a����5걙��e����,�ߓ�ƞa�F0~]~3zK���H���j}�_�1�O�[�'�ar��[�Q���QmU�3]�X*�_������a���Mݢ<���)S����jXXa�q!�v��٧h��00��Kkc�t�!���.T�s!�Q���%�������@-��Y�I��!�R�� �74(h����s��9����:�A6����kG���q�n������ZԤ,T6#.��$�RY��5�8��p%�:Z��v����c�9Z��<hV�4@����qduB��/b� :԰�ӱ}���El�PY����F���K���y�p�c˔1�-���2���->:�]1��&�j�l����#���ƿ,�fT�X���C�QՋe�{ ~tщL&����h�â@N(�nLT�V����4'�1|�{��(�:_��y���A�˖���Q�*�u"w�؀E^+[���H~�޼i:�!�7Cz2�n �EF�8x����%���&ID�`��Ln�󰉰���DU��E5��E�yZF>�d�u=��J� @2��D�tn��[��g��{�����TC����	@�]_��B� ��FFM��%{���<<��������\1�ZS8�?���|.[L�C>�dμ3���up���2��ṣ��V�Lu fy��-g=w�_yEŢh�ݥ�@���D���O2�/�A�ņ���p�ߕ	%WU�@L!芎
�BдmP��v�Bs��V�)z�Z���Ӕ?Y���� �n�+I�A�P@l���w��fIl-��yD�Z&z��pˈ���^a��%�;�����h,Lj>GE�F߆�1��ja�������{6�]��;eG����V��t��θ�J=����B2��_�L^�=o��7d�����J�=���Tc�	
�m�3*Ng!�����Z���\�Í��sKZQ���ȭvm�M�OE�Y�_/J;��aYM�V���h"�����F���(��+�X��5)E���9��T�WÅ��y-�1X�Tg��Ph'������;�7��L������*j(1�n�ƙ�(b�[c#�I6/]![�g���ES����Z�:�mB�Y?�mj�4�v$^�.��>|H��;	�e�etC\m�������CN�K��M%i�U��>�SLl�# �Ԗ�)|;t�u��vba�~Мp�q�E�P`�����O@�m]�\y(��h�yMÝ�ߴ5|���`=YK$���j���XG�Wn\���X9%��}0\V�#r��j��
��L��S�?Z��L�N;��s6��l�G�㿤�R�L�%%�ȉl�R�
�"_I-=f[�b;�=7�{h�";�!����!���_��ƻ^o<C����X�I�z�$�:��:O���78W��f�;¹L����n]'�y&L�ɡ��g���g�ˁ�U�O�C��.-{����륊��!'�r���\?��DC�uOȶ���y�XgҒ�5�(d�xJu% �Z���N��CSW}�#Z��WX"��t��� �3oR�)<���p�b�B�-��s�:$��bMS�̍~V����ө���.;@J��/�{^���{G��Mɀ1I+����$�����P�N�P�j]�|�W�r��$S���x��e)�]���q��Z�C�����!ֲ���?ODEOȸ<�*�u��?��0�Pg��!�۹o%�D���"hP��s�'��;�y۽'�dg�3hi����0I�n�-����&��B6��J��Hu�ߠK-�'���+���=�˘����	�2Օu6|�[��r��
�C&���nOě��W���Hzi(x�8�욇�1P&z��f9�f�rm���J"k'i���^����T:N|)����D������]n�ƹE�B=�������I������ڤ�+h������������Z��b�=x2���*��qi%��`Gs�<��L��i#w�����Qq���0:(]�5'n��?D��Hb.%Z�n�-6��y��J�,<�f-���Zjb،����Ȼ�`C��@��Je\�$��h,��.(�@��`��Tj|��g\�C�������,L�A{���.�5 V�e�&W�g2�FH����m��"��yz�b6<1o������3w���)��h�1�*	�ffZBK�Gf�:C����N{5���� L��s!fqS4F7�*�<r�*��A�

a�<��N���":M�'�����.��Z���ˀ/��N܂X���\*�}θI�/��bfL,~w��pc&�:-��g��G'�����퀂G��.�l`gM����A�j#�n�|�-�Y����LD���F���t{BSJ h�]E �YRr��h�^����DL��ŭ����倖h�8&yW
1ma!���=��<��K�����:��s{�"���\F������y�%�g���:���%n���f��[�й� ��|t�e]�AO �C�HI2���,`�m���x�'Ê�޲I`�ۤU�$;�2�#�X��PI��g�r+���I�⭘
��>�0�ס�γ��y�}S���2�N�A=P���ݚ4x�",,
�X���L/Sس@E��sҔ�rC��X�;�;�t<��[���hg=�p�=%��+ҵ&J�J,���W��O��41N���� �o	��լ�0($|4zOe�{��Q�%�#;4w���?�'}=s/+�L����p�lG��&b�U�9�����Pȷ+����^��>9���Y����LYbБ�lv�O��8�nt����O��*����X�������N���6:��e��S�(��j�zS�7[�4�gP�&��}�(��E{���.��KƉ��9h�"!�������nF6��S�d�Ъ�e��O=)�A��9r'o��\�HE7*�[�@���q�N�+��^��"��{�][�W3�	2��f��� O3��3�2�
��R����~��."���<��йt�\�xǑ��*�dr!\ ���$��D��r$�����|�XP=�s�ʙ=oG����ʪ��ͳ�h���C��w>����a�L[ɖ�f��7�@<�:��Gb��@)��صZCx�
�6��"�e5z�Z���f��;�J���ʱ�V�S��C�o�������y�j�\��}.R�Qz��QK��{���򐏜"(����X�X�Z���AvSn�����Z��z8�ܰ��úe��/Ϳ��@�*�$K$�e�^��A?�zuIhw�'[3HLT@��>8B�5s��~�u.g��E�<�h��vJ�5����w�p�T���5��nX��th�\xv�%)��}��E|ht@��X���B���a%���a��5HRx_D��W���
���?X�F?p?ԅsun'�D'W)��I�_�l���W}�wZ��=e�l�����6W���Xh�b��Af�U�����NΧ�$��و6n���-��+�~P�^�K �.�U���r����i��!?d�vW�����q��A@��ϝ.DPU�_"hF���i�w�E<�S;��tA$����_w��}6"eL҄u ���7�b�a�c�����#�X��kCAh	�0-�������H���!��fc��!}�L�}�F�
R6#��ts]�R�r�<�� �jp��z*���b���jD��E�\z0{_ ��M��~��yTx��ܖX�f�7�U�x�="�ec��P�Y���sZZ���(��R���� )����@����VW��%Z@/-�����t?vf�|2�D蠐	�oP���	�\��� ����&�����k��Q+�]d�>��t���/9���uHH��A�����'�+������3����c4������alF8���*D���S�^�;�FA�>}H pC�>/��u+��~�40�����faG0����ҍ�A/i��F2 ϶�m�hM����&��ꟳ�:�Y�v:SkYTZ̓��f����Ge�<�{�	2�R��D�l���궹�g���˫�_o����S�P���o�P�I`�8\zцeg.�]�d�������HӋ�C���窵pV� �Wvz�`�M����D�{���I�(�8L\,�5@8�{rIأ��fϔ�
�zz%c�+ P�E���;�:P�����Ȧ��O�+�4L��5p���L,��ռ.~مjnJ�m�1���K
�<,<v����/�6�|���a���VO�I���B<�D��;5��yq�������G҅L�p���)&�E�*��_��fA��k��ޅ#�װ?���w����!�<���G�6��S*�	�<օ3��-�i�,>=�o'η�Q�rWE1�ƅ%�Q�{}US�x���Ǽ��������}�_UЇ꟨z���Z�h<JO%oa���#1�y��� A��;���nW^�}i�j�B@ȍ��e��b���
��1�L�#$�ļ�������:@&B�Rc�����W@�'�㷊P6�E�|z���o�o�4P��p�(�%��lݏ��j/��a��X)r5��١%����7�j ��}�g��ޤB��TC�a6��H�O�਒G�}/U[5��iز&���Q�O�|�"0g����M��͏��xۈ�}	|��ы���k��1a��p�gu�s�MU�����!F׫�Jhn�#��zA�b�"�Ͻ����Լ �g���`g����-��m�x��U�qs�Y���e�_$��1�K���n���1Ja�ǌ�"�Q��ɼ�0I�e�C����S�ۯmHו��!z��_Q�"��~YLi�9ܯx��U���!��V4���>\����cO}7�Ҙ��i8�,��L�b!��q!X�F�Y���o\(q���/K��;ϜN8,��x���`��^��*��Qa���#�6��v�[Gfq��:�p"�e���P����7[�x�	�ܼ K�'�L>�,�I���+��!w��\ ��6�᜛k+:^�\	��yo{�!���F��dˠ�~���7�19��n\^�����ބ�R}���Y3�|Q�{�UY�^ �s������K����m����jx�,�{-J�O,Q��ǂ������W�F�D�r-��Z�s��BS��沼|`���ב�_`�&/Fq�'�Ip��JO9f5��Sw����O�ל��gJ�;�Gɓi��I��9O7�J	�7��4�ՎJ5�2�1t�֝@�[�d����lp�髈˓a|
�)�����J�`��1]Δ�mcG��_5W��Ւ�Q;����8���Ֆ�'e�Q��~��^d���O#��O��{�b��?CW�V�L��_lYG�u�'�6�̍c��y'��DZ�38��&x��Ȏ[��z⻳Y����r�`��{kn������Тr�����e����8ϧ���/,�cuZ���l?6�2e����xD诙�Ig{�[�6	ևK1Ɲ����J��Č��H�Rɳ^�����p���,[�����z�_�z����;Q=s�xn�fO�3* �Y[C�4U�0jI:�DC �_r�<4���k7PosG�7(o�jR���_��[a),
�H?�H�r�1zQ�=Br9�̙ .r�t�FL�v �M$��W��A=1^�ݏ(~q���&�㽟:B�ѿ���5��$��rA��B��d�%�B���3�H<ήF��A�ۭ��p�T�y�m����O<�*" 1�apȕ(0(y�0��J�O����Lw/R�P[�ଞ%͝��L�� =���e��g�<m[�Y<I��v��8�/�j�ed�i��yT1&N�K��(�q���(*!z�5��F��?m�����5%>D�aLr�r-7?DNC���~��P�O�O\��j���T©����{<�d����Mhq�L�|�.C:��w"�� �>�8���-��R��D&ԡ��e��$�
�2{���'�mR�z��ł�p��QO�/�"���Z�3���r�Bg[�0K��4A1��bk_�C��DUB,�忶四չb��M��3�.�Y���3�Il�H,t��"�iZw��.��P��-�� �e�h$����Q�i3����r���J.%n5&�m$��
f��<MkO!��-y�4������hn5���ȫ»e���D(fI�� �߿A���z��;�Y�0r������G͡M��J�`R��u����Җ��i�^��,2�~�:��[��dun��$:�5!n��	�e�3k�&H��Auþn��al}3q�KPI�oܵ6:�N%�a��z[%���	d�	ё�RO�77�C�w����<�!�CIkd��`�(���Yš�=���~r S�|��Ж��ӳ|ð3t��2�!��-�z�j/)���AD!�:�� ��}�D�(O�c%�$��J(�5��#Ǖ^C%D��P��Q�y��R��F�<�6Yek���w�[祘�6��������H 4Sb?����ד�Xg���I��;ﾖVI�9���*�}��1�+b�FUNf�p>�)I> �n��K��8
/��ޘ�F�ӊ�ٵ��4~O��pU]l�1�W���!�O\z�+ȦW|8�©zK�'���
�ӰU���7>U��H�4f�=0��F��a۰�'g�"�Fg'i9P��f�R?�ůg��J^�����������QCG��Q��}��,g�7;��6[	�%���F6k�������%VKni�Hْ�`I󬷍M���f�G��fR��l�a��b�R"�į܁���h�!��m����!�i,�U�cwI�Vww�
�_Q�Y?vM����`�K�=
҉�r
�l���ϣĖ��C�S�׏�\�(�A�F~ .�;�?�Pr���i�yw��Ԧ�]��Y�:��sn��5�$
E+�ǡܥ�{#4�]��s�
�A59�֩.�2��*dO *d�>�ʟ.&�"��6�p~���)9�Plh�3�-i�P�(���KZX����&�n`[�3�q����a5����I�s��}?�vU�iX�Z#����^��LN�O
q��}��~�{�Kʐ)��� ���Hޣ�I�KO��q��u�q.eըet�Eb����^>�hW�7V�;A&����v	q�F�2yǤ\�R�_4@�����>��K&�
Eڸ�v��"���IjT���|�A�KY�� e����]/�	�pz���RZQ����+��.dr��䨭h/�U����sB;.w�8(�c���U�C˅��Ի�Z
�Ĳ�@>�{�u���([ba���W�?��K>#mv�|~��\�2�bq[�y�'�}8Qȋgt�!��O'JjB؊s�����x��AQ˭ɐ�4�6+�,|�x�&�HGH�Ի ����H�`2�Y���p�8Jt˅HT�*4�u�LF�\�J��PΪ�4���ڙ��LNln��#�zJ9�����̢�)�x�i��1��?t����tǯ����e���hP_&��R���Yo�ʳ]¤2@Һ��M��7�H�P��ҭʌ���g�Y|�Q
��`��Πxʆ}����v�ϧw$	hv��}� "�U��;ڛ�����%D߉޷N�����{����V������T��d�$�߂�	��I*W���v�zC�w�����P0�~��Pf'�\�1lwA��p�.�b$���%��)\�3�:�f��B£1����ެ��/P/��eq"�}�<r���yD��5�M�G���K��BRM8>G�&i!���Q~�],o����Ik��ʯd	QB��V�'�{�Q �	�$�-�o/k*�=�$)l��L��&w�v[��4�E�V~�A�Qi���+˻��%�Bg-6+��������H��3�nMFLY��g��Fdl˚��%���r�o ��T�J����,/\�*!�0�8�|�@�J�V�܏��^'qoC��0����3oo�b�j0;�:tQ��L2��.���dk�0���a�H�����ƚ���5/����L|(����%��Uen8�����A��&{$aX��"�\[��"�����/[J.���*�z.�6+�>`�q;c� z��_�0�����F�D;�5It}s�H��qQC̷��Q�{r\���!:1�\����P*�YH��|{�8'o����'�yΩ���h+6�2uv��p[�������+�n�E�����Y+��y�	k���r���5SAV�N�%��&�� �Ѳ3fK#�}�������Ƭ�J�T��8&�<2�C�E΄���9�����V�0��ֻ���z���/� �J��V�2H�
M&�J<����>RZ�ZN/c�$�&�!��"�0lU�'s���4�N���S�VKk�E�@�Q������̂�!����o���6��*ԁ%��1�kҐoA��h��'BP��\.3y�q:����O�a��==	�����oغ���}{G8���$�I�i�4$��!O�U����k͹�_*=o�Z�j@��X�	�V�SA#���S�l�&�e�u,Q�����=;�Smt�~S��S^A
Z���b-�=[�����t8�wt�[�y�L����,m�`B�ހ�GO����M�U��8<%��Tt����3�.�e�r�{r��=&FZ��t���P��+F@^�ۥY#���=���8N�F���W���hv����	3�=_b��3�qB�u�_����O���5o}ݰ������L���C���p��L��	9R�b�����txѬx$�K�~ky�Z�=^Ҙ���d��ɣ�4�����4��2��D+:@�f��P-7�+���|��������!qS���D��v*��|Y�����ⴊ��Ux��$�u4�7P������	�̹���y {�`�O���ܿ�ճ���љb�g���nך>@���1n�C�|�ꁯ��R���&�����OTr�?�9�$a5�"�f�w�K����m�|��~����X�@���R��z��&*l�T;[`����LibQC"ڲ��p�?Y��Y�!
�����Uv	%���B`���a���˅E:�Bq/�;j1˽g�G��������%l}�a6ф5|ć b���zG�������<=��f:j��^��!�� Є���)����ߺ�}P�=.&� �y��O�a���\+?T":�D����o_S����!����5�w�J�Lm�e_5��vVE��`��廖=�(�&�bI�4��8b?g�ݪ�@f��g8��pz���@fُ ����G�KU��$��³<]
�i�
��%��M�+@	�;92fQq\�����l�T���K=d�����_���ȇI��Ƹ�>�^�n�	���$N���D�D�U���c0�Z9g��(�J`�:�dУ�F����C[H�ޑ�e�����d�P��v0���Ox��m"-���X�����:��t��V~�o��%X�Q�ϣ�
� �Ve����T��wD%	��]�u���ѐ���[q�2����,�;�A�-�k���VaV��mF��kS��+�tr�e~�ԏ�$� Ywl��A�
ٶ���rz�v6	C���{e��Y��ھ��v��l*i�xD'����;W�+ {�R	��G���:����f��#�٫�����ý���2�B��R��c��Wu��d<�E��5+�֦�)8�� V*od	�qY���CfB�������*�pY���R�!0h3�d'�lk5�\Pժ����v����NME��U.s�$��'rY��e��>n4��/̇�o���1���D1S�.2RM_iƣ�C��ֿ<M
�T2):{���湀<i�m!��N�}����4��,ll�!�	����z�(����b%(��z1a �,^��S��(�9�jm`��W�� ��'!�s���;�$�������s� �
��S�ɈRr��% �cUP;3%?�##3	�6���Gp��}9��);y-�^_�^�\��y��^'T�qH�����}��������u��%U]���A�U�LL�Nd�;�3ʵ�Bd�e,�S�
�:i����M�>���*�C�_}����}����yX���q��2��T���wc��V�&:���~��<
�#�����.̳:GY���O�Ob��]�� ��3%�UZ;IFy���}5Fe�#��~�:擹}Ψm������t�'��Ql_J�C�������f +��§"��x�@�lv�k]iQ��d����Ft��&y��JA��>� �k�(��g�� '-���sSʇ̂D��י��(�1Pۃ�����'���p�<c�e05Cp�=[�N�9J�1k�$e`@8(�(��X�>p(�
��	iI��\'�������YD�BS	�r{�Ps:�wD ��+M>��/ԨzG8]�O�֥�.��z��;�p0i��}OdJ�b�l82�c�r�����|�_1���C#۟cB�~7�h�Qz���V&Y'��|��gp��/�:��f�7�x��EZ�c+v�ap3�X���ow(��a�@������7�Uû\d�'p��:�0�FR�+m�w�,���$y��޿��������d���5�Ѝ��x���L�Rw=)牛�W�C�ͽ�N؃(�gݷQ̊Zܓ��y�O��ף*ĵ�J���%jt.L�Ex�G����||}�n6F�t�(�}�Z^nC��7�ʸ)���~w!V
~q���r!n���r'3/!���(�WQK6�%=}NŁ=Ϣ|O�jχ��D*Sc�R�k5��|���U�ף9[u����R8"����>+$2v�_x�k�ЧJT+v��xr���'����]O����W%�3FXU]!a[�ltb1�孎{q+mk�L�>�ξ�����C�(
*PH�ķ�3�"�J�^�s��JB=�~*a��Gh͋�S�Y�e*�q� �Iu�y.��`���x�6�ܰ�`�j��!����A��B+�#OߟBtu����	dBrn�[F�Ds�ϑ^�؛ H*j���I�)_��L4���W�@�����R��>��v�0(��[7;-#W�-�4��X��\��:��#��6оBL�I��z�7���O�V����2e�`y <<�AW���l��Ea��9�hoy��&2ݕ0�g6����(|Ԯ�����V��!ȅt��#Q���un/�N���qc�೤V&�@Hd���n�~:���_Cp5�a�W�j�A�/��kb��D+x�q\������'%�I��������K��Q�f�����B3�_�����U�=�� �3H���.��4�v��E|c<�]�O�K�Y�C�r]`��g��6�lj���;���D�&�/ ��=�X��.�C����n]b���@�E9Z�TE�&���G�$��@2���+���M=�=��<��$�	1�6��6E��Vc���M�
m���&���c�kW����IU'f��3���E0�l�H�g0�|�<[w&f���w�@ �Maߚc!�E����S���66�,b&�4H��C�ggPk�dA5��'��'<���˙��YiŶ?z��^c ��il��Yr�_����D1���c;���C���R�T��i\z&w`&��ՏZ�xR�� ��b��,�PY "�,}��yֺ�C��>F��%]�g(fkh�B�.k8���X���y����0Ԥ߽C癙�>��}g���
E�-r�yr�ch6D��b��r�u���[7���pKAg�2���v���(l�E����J�ٲ���fxJ׶Sa�ڵ��::�wNhZ��O��T���pi��:��#2�C�+���̘��n�\@Ǉ�Lzzߎ�E�Fq�(�����}�b�s1����L_�,ы��Zp�1>6���`��c�]���������C�;��w�Yۿ&E�B�Rdn�3����V���f�ѥ3O��t��r:��M.[U�D��ܵr���!��b�G Y<D�,�.��pƔW�q�	�������/� TG��P-%����Pi�R�����Q�ZF��	�-�-Ir�z��ˎ~��6�+���D���^mI!U8׆���T�yƏ�
������U�� ��S��E��FS/S-4��|��,Ff	�6��z��V/�2�,���	~2�1���e�Yt����4Sӱ����ۡ�eP��9y�-ɠ����&�M��˛�mc�'-��4?�=&ު#��ڜ+do@3�>��}xv�sU%��~iL;ߡOV�Mn� ��k�����|�[�'a,$��j����Q��IDo��h����P`�eR�~��1��p��8�����`��ech#�3轥�6&��ibE�6<�EZ�322]>c���n�k�Mm��i���6F�
�g]~����6���/��ɾcS��{��Lꯋ(�n�����f���+e��ղ6=�(��e [�H��7�|w�;��tl`Q�2Fw�pџ�4�~��k�}�:��N��NYNXT��QVm�:�%1�Y����SZ'�+�>�ʙ�t��3E(]2��B�^:��tt��y%��9Ou���ؕDN~D:Em�r�������ك���;�r})^�Wr-Bi|�C?E(�]\I�g=!9\�-��=�hN�:*s�V�2_���j��e ����ӈUv�ٕ�� ��[����<$��C�`h6�2}�I�/�-)�HT�8�rsר��Me�������;n5�˿�a!����x�@SLຆ`;M��D"�eT�b%׮i���:-�(�Y���Z�V�����5r�ˑ2-�M���U	r����ĩD��y	����4��q�g%���ܦ:�>S���E>k%���]o�N�ד�g�r �;ƬR�H����܇g�A�7r�*'T�L;N��Z!����g��	��� �\��ƴ�]%�~��4-�zqmF\���A�7䣟֨����-���?�N�E����Cs:�������Fp
���߯�m�kP�D2J���8՟B�: �t0j�3����2��,�/@F�Y.B�y��'�'��ʦ��;��¾p�z������a�p������H������!��$)�g��A0=��3bQ!,���xJX��E&-/���,n�MN���0C�%L���h��h'3?FUK��;�����<�J�Jx],s�� ���k�Y�O>�/W���\�w�� �>,'�rW ����M9��V�<cI��^�B��#`v�"��Hk�X�Ȩկ9a)٣��^Q���,���"�$_����:t��榬\�?	���Ҵ�1w��[�|����s�e?ou��"�y���yE�Z�A
�U�A6�%�:	���P ��՘.�VS)4^Tg�'Wm9Y�x���6���y��be#�����{���S`U�_ju��*a"0LZy("��θ0y�"]��P�ȫ�#Pً:��[����5��센� ��-�C�T�@qĦ���[Ƃ.@?g^�ӋY���K���#�5ta�{y���[�jE޷���/A�A��+e�SP�g7��r�;�׋AߺՄlSZ�%zD���+���R�\�2����e�q+A�m����������5�tY�����"=��b��大o
�x��2�xo��ʊ��'D�BTP�����S���E�-[7X�~�	�@ �B���Uu`X�#�#X��?4�Q���K!wDТ���P/v� 2�QM�U���9�0�N�!r����4<I�O�R�c�f�v�K��7�{���lF�L�e@Ϲ:�<3r�C�KOE����`�!<��z�n�|���-���Dȼ��Y{����k{�=q-�lsV�f H�s��+`2[y6T[b��F=H��q\?�
$Ï�Q{:{�S �lk�ko�PW!�Tq����kB�@�5�_M7�H���+��R��7'���$�p|�:���s�kl�=�ɰN:}�OW�E��7���%'��:p7� d!+��[�z�xR�P�]M-�gm󧵵��k4�*����̗%Vo��qb�e8��b�͵���f�r%���\���C4�Q���1�y]-�0{��������"�"*a�"�/�s0b�07g���
�niM{���(�A���HX}mY�>����g�%מּ�'�<@��lV@jc�zѕ�nymݎw����|�Qa����$t�}G�b�����j��wi8\�~9�h{�i�-Q�,}���G�פ�t�t��Ю�C�������qxRQ:�� (�p���;K����J�(\��w񕡳��k���6�7#?����ا��N�E��-�R��v�+d̢l˨�x��������:*^ X�U�ڪl@�;'׸	]KV](#z�ѪT<d�Dّ�4wdw�J��U?�;J#��������4�H��
Ń3��89(�9�D^�:���������[b9.#�X̀w�����`?Q�T�	��U�7*���O�_D��@//7�W0���1Y�H��!d�[��l���r�	�Q~3xr)x{a;�`�ԛ^��-82#�y{+K�
o�B�݈e�Pbr�C���I�K���|�$j5�K�_�u?�;~%�-�;%�����@b�#��s[�q���N���K/⌾-j_X�σܣ�,2�Q��(x�$+�D����G5m>Ȫ�� ��@��B� M7��@q�p��Xj��x1#�pa�a?,G���|��#�e�΋�1ep�>���n9~��Z�Oqq/G��Cκ��;$�`�4b�&9�C�7hl�ި���7֎��<��q>>�`_��*�ڃ6���.|�UGyc^��g[Jv6�z�!��_v6�n�&O�ǡ~?s	��oY�b
��զSRA}��x�B#�ꃥC�i��3�#���rs�	.��Kw?[��e��wpa��W�F��_X��]#�ΰ4(^jy�5H�� �P��T��p�5���6g��g6@3E���	f�E�Q�"��2m�#T��?G���ѫ����"X���L�2 �P���6�傿�AԅP��1�Ć���k�>(�:�%�t��h�8;T�-GXC�b�ܱl���{� �����W�
AQ9#�/�ѫ���x�D��X�k9=���xD,��ٞ���^ �#�N1	�D��7h.=�ieb�`��9K�@��lNu_��<^��D���@L��MC��8����S$�r<9��<:��T��Q
���sa�V�;��[��[�J?#A�%���V�際@7�i>�6(բ�;�/�Q�Ko�A��aA�j,-C�|_�=�;D�~��4�V�0�g�kP⋐iB��	j�bFz�O˗<B�5�i�Q�����{50�,fS)9��E��E|����n����Mm�T|�ve��6גK���(�����]7��1��/H��v�2�>`'���t!�[i�r�Ŀu6\��O��,,D5���
��E�x+0��x��7I7�L!�`-D������M�N�:%�� WZ{�,�(kQi��^9/L�5I��.���A=�]B4 ���E��I�O�W�T�q[�T5[_OOO;(LA�a��+���+�����i2�b�;���R��a%��nn ����R|y\!�bs-A�=�B.����o��X�]&d�\֞��ȓN}Ҳ��
��1�|��NtK1����uM(6B��<�A�'��l�%�c�l��#�iQRۜ�yx����wk�HiH����+%��P�\+)^���j�h�f�E�u�ʚ�8���[��g&i4���fM� \�˝u���R��\}��>��2�ӕ;.b�k?qH����b\/*� �)ߟ��#�L���X�����$�Jo�G��6Y;��Hb�*D4_�VB�}Q�Qk�0��9Z#T�c9���`�����k�(d��	�a�akA�f����y������J��8�W��2<�M׫bb��8���s:uh�n��@n�	�l.y4��WP���:d�$������W����K1
��+�R�JtR�EF�2(T�?e��7.̡DT�.���-��E7���#��\�s��-�lh����sM��Br�R�_���&�>-�u�T�Ϲ��\z�3�VYrZ3$�
����S ��L�:β�0e[�t�y\��1����3&��	�#��[��2m8+�9�zY"6�J����yI[�o��ϱjs���d�6����Y�8w��a��\H�\�V����W����5��g���"����M��]�_���'�����㤼�<��d������C��͋H�|��v���͊a� Ă4��:yF3,��������x��|e�*ln�(�t?�d����?�������13x*Q��=߲�F�J�i�-��	���}9^ܟ��]�&^��M6��f��X�S�3���NR�G�C4��V[��D�B�a��#�7��6�`���@3m�FF�w�aG����չj�ݮ��r]����a��IW��|�DI)�/F	�k|�rn�&����`�'���9�ٹ�~	��b�!�n�0k��ۥ�I':��}�7�Sy֣u�@��4�b��4���^�4��U"�D(l����^�x�i�N��Nr�x���Nq��ܯ�N����V?�,9Z:�c&�Y�]�/����:��?�ct�mSZ��0�,L�����S������<2���S� �M��:0ng8|v��HBV 4i�~�z�K������Vp�����
����C�늿�s��}�X9���	%�i�r�kH�̓ޟ2�?�%��,��fFA��N�}5��<��6�x�U������_c(58�Dv�:�i�ܬ�F�#��x�[�����_�O�-���T�JZ�ܧ}����I�����]�	
[f�������i �Y���3p����d�=�$^�Jj�y����/��sz�Bp�����Ca6Q)�phUϟ^f!^u3C��i"�Ⱦ�
���ʤ��TL�_���*�:q�`=�[i��/ffj<����_��*���»K;��u/U����C���� �n������M����+j�3ҢB�m���,�����ѫ=~,K��T����A	���$ky�GBh~����t����*K$����M�C x*����a���5(��|�C2�'A�Լ	Sw��.���i��;h�f�>�3ً�/fЬ�`�bF�u*�B�iDHD�t��TC��
nM�s�p��Ѳ>�Ӣ�/c�kJ)����oш���T<�t��W�;�s嘆��S�c�q{�qe��Ў� Ɣ�����$pe�aD�c��d=AXPE��n���z���]��ʐ�ُ�{��O��7�D/��u� �]MlK-�L���3p$�P�N�:�M1�0�"����]��<C2�T���v۪�U�H�%��s��O�TԤ�&�K1��RY����d_���q|^��]�Ж���E����y	i��j�����Ze@����1zoS�&�V�C���Q@_*L���[����0l�`�9q{��%SU&Ѱ�FU'A�� �Mpf^��crNl6+j���,&�_V��VyC��������q)b˛��W��'ul�/$)Q>�]����4)��������[���C뙀m�p�[�@�����a��RBC������!0(�5�A��K{����M�xY���1f��"��i聁�0�ɔ�P����[/�En�P���~�Q�3a��5��G�Q��L{\O�oz,�r���m	%]d,S47&s����!�o��'I9�Uj��9��
>�EeΣL*E����I@��4��1�����د�Xx��>�A�Q�-���.�n���<�Y#L�"Q���F�)jm����]������Q�F� ���Ul�o�t�f7b�	X�I����6�G[��&H�y�1��+fW�@"����*لd�����7�@Tz6�G��;v��T�.�S3BV�ܬj���A'�[��*�㷱�#�����եWC����g�v�Z�lIѪ&����Vǌ�Y�8�K#������u)DXHH
����DrI�@�Q����h��c�P��86(�UD�߻����ð0Ϛ��&QQH�bL#�϶"�1C�t�3�°"�^�Y�!�����&$؊��NvrL���9&v�	���}w�w�L���y�y���׎s���N��n�R�z��nCGL(�2��V��%�p��(�7g%��	�3�p�X���6�vD\�¬�s!�RIw �/���l	�2���W�����ˑ��ٽ\t��k�k��l���q}��"�<|3�q��rU��`�i�9�����v�ەU��c<�ɞ���&1��B�%�2��e�[r|�t-��hLE����au�� ��8�����q7Fw���j�,����<pN9����y'���ܹ��_`G�	K8ʴ�C�2�z�栕��~����ċ	Nr5���fv�1,20��2&�[|ibY�;ߚ�R���-���h3m��gⶮ4��g�0@8����� "��n�2v"w'
���a*㻪��nhm
�L�HPC�s�P5pC�f~h��h�i>�0R�v��]Α���P��att�D)���8��1ԑ1ϮQ���:�66�xi�T�d�C���V�����4A*�|mW/���z��k)�E�*��C�v����A��Z��x��+S�G9�=�m����ˑ�>��/<�	eK
a���|�7e��قT�}�%?��a?e��,�j��m�@oG@��N�4)H�=ވvl��4�x�>�̟���t��S8�ﲩܛ,4���1�mz~�����I��j�9��V�{���Em���u����V��S�9��$�x^+T���*��	vX�@�e�%�+�݊/:q�X[Ik[�1,ݏ=r��5��͆�q��u����]+9K	nGe*�֍����ٟ��|���C��%I��Q���v��Unl���U�����V������s���A�:�%;��E�v�*R^��@A\�~	����2�󌰢��E�r�TX�zs^L~U�3-��'�y��~���Y��D���%���l�c�i3�wҢܻ�k`��VԘ�,8ؗ���$�O��uP�F�Q���P����� }�'EMk�4��N�e��m?���6���΃��=&4���9'�-�u*)1��aI`��m���t�-��4��R%�8T1��QRe�50���������x���/��c�Ǯ-7�S�TS��̍\��M�A�$�_[o�	]H����$�.nC m�f}exO�����- x.j�
��5Ȍ��;�r��I|��|�§�i����n,��U:�z���ăz�?��}V*�Z�>N���+����	4�sW�RS|�D�8����Ԭ�m���@|����Ժu���TsN���O.�.�S�V����S%z4��m0�'�}<m�֪��\�f����%�T���2�*���?��B���U$<���NI�fK(y%->���2��C7kT�l�@��%�{ҭ���ѽ�.�j��BճRI�)V0�~���F��)s	��o���'�<dM���Ǥ��4������G�	�*�"����ԅ�+Li+)XN�6��L��m�F��RX�c�e��# 3��[�^Q���%���֒�������_�d[���_2��U���W*�L��}�./��� � �7|沊��/{�zC�{����P��@0&M�=[��
��J���o��` Y���Z�[�,�iU��蜧~�*?�As^��f[�)���d�}Wv��϶���'�Pt�(b��9���++p �ĝ�zx��d�TR�)d�z��ƕs��#�q�T��+ g���i"�2��*0�6��,�Q5�Z���%_�����Z����]�=w���k���F0�1�? ��`��0�Q�����~��(f��t�١6��Ŕ��Gyw�� �}�D~�K�b+�؀w����ɒ�-� ��H�ZpS�%ƿ�.t��J�4�׎�ֶ�mV�IJ3��q�.�����9��ʇ�����ѷ!o�����a�;��]���p\_�[K:a	T!��^C�w�,STU	�]S��"B��yף�:D�e�N��vҜ`�o8�l����F;������%���qRQY�e�M/ǋ�)'��kɕhi&q����t�M*�Nm�j�4�bF��,9 �̻8k��o�֛�&��L� ��R�C�[WtL86@4������`BA�N�b�m������dȫ�u��������wO�����D>|��#̶0�%~��4̈́6��7v	�=����* t��l����v�Fs3���/���T9��z�Ғ��|h��g&��g��j����)
�"�HJefi��1�Q��!���zy�����R�I�[;#US�#'Wb�a�ײ�^��Ѷ1Z�B����pŒ|&A'�65��vº_�{\�""�w{[Z����Ɂ�����B�2m,���uQ�T�iFԻ$<HD���uaqi��f�!_?��\���A󱃽V�{�Ī���W�A薀��$:����9\r�Q/ھ7���^?�։�����2�Av��=J
�9<��c�h�Vm����j�n�*��t��\�͈���D��P�2��a��k�6�e�J�O���2o��D��U���1;�����G�t޾k�1�aK_�Z�b:����&��Ȁ�C�"�e3|�i��q=QS����?}0"���:y$R��sly�^-�T2(mG�S�Ty�����-מ���W,7ycCl�J^�� ���t��G��[t��iZ�w9�|�P�m%4\I�o�����}�iU�o��tRv3�	�*xܸ�<���L'L�>�}�t�h��ܓPY�
�N+�o���