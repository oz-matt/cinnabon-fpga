��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]k�j*�Q��~�=�0z����o<���_TC?�];iW��M������O���R�$�lIlqֿT����N�B���Wg��i�ٝ#ei-�#�D�ዣ�I��n��Ώ!Hg7��@���ֿE�Yy@�����ɰ�W�t���<ņ;P�J�R��J}�f/�	En-Ԇ �c�}�g>���C�&Y��ȹ���d7���F�<DK�1��īa��7���y�s~�[��d��"��5�f 1�?w눁��]�"��2��f<ى�ʳ�+��-�퇌��rSԎ�������@��Zx|^���E��_Dj�r�m6��n�7���I�" "Դ�V� N�k�dlO,4^��)���+e�F́�Q���iOH�Z��`�ٮXd|�+����u�q%��<7?'�c4��x	̶�$��۲e�e�;:Ol!�M�:�>�+
r�3%��'��?z����!<Q��I��4S��4xM]� �n=��reB���>a��>����E�=��8ȫ}G�����ׄ��dgC˥� əT�O:?��kq�]���p�X��tڊ�A�	Y����+M����:3��D�_�.�Q͌,�zQ�\�a���Q,�Jp7#�z���q8���N7���)�x�Z�aF���g~��%i�{��$.e����ȕȇ��+-��?��vx�R?���X���e�G�5{��/��
_ž�lկz�sĠ
M���Gɻp�;��rT����i*�g��{�n�+_d ��iX���-�Nn���-��cĭK��n�O����o2oȺQ�F�9��ѕ"��\�dE�q��lƻY$�(b�a�٥e�1h����m�#V�¥%
n{TL�A�H��ڨ�Ti��f�Q�<����b�~�� �Ƴ���d�V/ǘ#S��`[�\�E�tǹ�e�AקG�/ ��~�+�G�FO��"L��V�q}�4<��G� ���Ka�з�T�ɴ�%��=<�@���g��^rJ��¡���Q��$
i���~[T�H���yʶ��d�Z�e�څ7o'➗�8�-K]�6�?SNA��z1W�M[����0�Zj*����l����'�EW��!���Vica�PM�I��k/����b���\=R�0�C���haQ��3��4y�N5�ڿ�$N{�I}�"���0/oB���|�&U{B�� �o�07t.dF=L{�`�?����TD�+�J��S�� ��o�N�`��n'HwƄ2�'�\}�N�.x��N��~��q9�"�+=��,��v�)x��f�iN&f�l�q�"[I7��~�@�z�]�����`�Z���8Q�i�7�|���c4∿���w+�0�n��i�:}"VX�ZZ�BbBik��5c�y9����oE���r�"V�wr?�gy<�&>��1��4C(1�������x;��4�؞�F^1�Pũ���}����;6�
G�~���R_��+eM߸���K��^G�������TnK1��!A����������[����V�<�������@�e�KY��<��������1����Ϧ�����4��:7}����~�`ګ�/F��'�F	Fv��1wG�k����͋��]9�l�������2����ă�'ހX9��|Yš�0b� ��|�Ops%�̩��q͜���a��S(�1���AB3�(�	Dӡa2�30����`�D:7��.�p��H�  ���d.4�-�lܣv�5��U�F��Q}T^r=�綔.�R��1�_�B,��:��VVt���=L�_;��X�m�H�81����3O�}����J�-d���o��s�3�#���!��,6�3;�h�:���I���`4]��A�,7[��C��8�hB�
��ս�бj��b�u��K�:�}C����?�~�@tp�Z}U�B5(�q�|w�)IV�'NrbhS/᠉��Gu6��l���e��t��
��&��؏���~%���D��3�U���[�?�(������r��MzG�o��pF��q�J#L��	}w2w�R����D��x�ҵ���ט��[��:``����vG��r�Ml����d=�?��v^xҊ��6���ִ��G5wmWF/
�^ ��Q��K:�ɣH�ȯͪ@o�x�г���� gښK���BX�7��#�4z������K�%��[�'����ԁ7p��s1�ѽ!)�޻X.�1$יn$�������m���̗yT��_� �"qH)�;�ث����l*��%kU�a�����X��{���{�5���R����a�ݬh�5�����/���'GHy��(��ǿe��xI�0z�Qs�a��3�6��Q�k��\�U��lҽ�+^"S����~�TiU���wN�#�P�d���&�՛T�ś��U%HQ����0V��e���X �W�Vc��oP�}'c'����1�F�l_��F<>qPpzÄ��C눏�&e�V,V��*��X�2�䒋n����RHD�y.�/�u����y�0�#჋��U�n`{/��_?�zR����6[���CO�IA��-��O�P	�#�3b���[��J8�j��/�0�����W�+
��t!P��:�(6������Y���b0�f@�b���m+v�3�,V�v`��8�-�ϐ|�T�~An<������R��.���3�{�ظj��0&Xم瘫ng^�:��cĺ��fL���6�cF�'5C�A��X�Wg�ʎ�Gf�j��ȯeO�]qh�Ȩ��\���2y�}�3�����Ď�h�aJ���O�.�G�-Q4S�j�"�$������
�% (ؑ�OG���h������!f�x�G�a�@�AFP���i;k�K�v�?m���t�l�Ӎ��p��A��@6� ����m��� r	�,����;p�,o���l�05R��JҸ8]�5��(�,
���8�3���q��yw3<����G���zj37^�W�����k���~Z�������ߖ���=�)e(k��^LW`��y&�.�;��U]I�Zo��Ӗ!���
�= wNd��")�c��ׄ��(��t'�_��8ϙ��;D|���!<��)�%<{�Sb�ߟ��Ӟ	�%n,(���e��1'�>Ou.0��r���X+i�J���i��ю�G���y��@`
��r��^��=����)c$�{ˊ��aRy��GM�~x�w�5��ۮ`S������SW�W@g0�X$�
F��wzs~�@6ه���t�[�Q��f�qq�*�6�FTi�N
�y�U����MO%O��$��;7���,nnά�l�s~�\����h;p�4|��o�!�a[�:ʗ���(���'�ho4qڜ��kT-�[��U��C��o���W|�QE�r��6 �4
 tX��s3̼46������M�<Ξ�vV��͝���m�}8	����
�ۈ��.�B�N�G2ڊC&pX�%�/ѡ>gֶ8�V�\�bCy&:��Dv�P�*�:}�-�vP�+� K��M��k��62���}�#3+��돁
欅`�4��{4�6�/ps�����&����6�,ߖ��T�Ԣ4 � �q�k��%h�l&�p*X?�����ߏ�N7S���1��âZ���Ӟ7!+���F�"/.$�}�E������ހ�������lk�'N�o-�d��缹ē�䓻W�&��+L�C�&�\�AJ�]�.�1?2�HjP�����i�N���N�J+��-�6)t�!�!r����e�qf33�������@�iM2���#���I]%2�ƕg��q@n-������&t�^��{��e[rL�D7�d\�������c@�k�a,c8+MZ��h��{�� �Ϛ1�e���+�y�-���	"7�G]La�_#��5����k8�`����J�k�h���) �}�P)�2�`�-]V�G!m!��!�^����c�G)ⶃ�:h�f�j�u:�U���������O�ǒ�#����
	U�}��deE�jA�Ȁ;ﴅ:�)��9S��.c�Hя�X�$��l��2��ʜ����q}d���&���Ů���ܼ.�x�M���LI,n�� �g�>?Ó.��y ]�h�R�nlɢ��u�s��,W��*�'-c��_�=���v�7$|&J̝���5�P�0i���F����*�c��+���l�(��W�f�e/Ǆ�����m�Oq-們����I��Kk�|?�}k휷��(�J2M᭸'Y��
�1�2�	HV/*-�0ș}�n�6����hd�m�lF��}YF�S�y34�ݡ����/���(��F�mkն�,��_V(G����_���pH��_µF�lۤ�k�y�-�^%����A�4Ѕ���O[������u��꿋�$�"���z���H��s`+��G��)��w��$V�:�G��	[�
l�2e���~ #�3oc��k��+�x'_�`FB�t	�f졿t�r��[M8�[Evv�õ���C�f�ziT1ʞf/H�ڭ��]4i.]<j`��!��/�S̿���Dj�d?:��K�B���hv�U�b��uw#�ڊ��T"J��	�T�RX������h5�'G���x�9����Ѻ�ؚ�䆧����4A�-Q�>�=��u��Y�[+1�s�Az�O�g1�dj�J%pN�w��ސzt(Z�:����i���_�wDbC�Фl�����碑KAC�T�+9��ܠ5�+�ϯ\�"�V����A����Lh�?ٲ�q0�*��ɤ���W��w�h���/�ę���0�r���N]I_|<g�29�}I�,�k�p�mX'��GIu*S���5���\��r�˲!"��J��q�|>;W5���%��$5-{��vie�R�|�_~��`��j��}AR���![�"�x���EޝA =�c��A[��;#��,�	3߼t�˫�#SF�����>���4Z�����Is�8���t�VZ���u�7�?��Փ�{�G���$K1�|9b��P_n-:���|�M8.�Xd�\;)���|2�$�N��D}�l�X���vw@�-7Է��ER\H�$�/YIi�jK/�j�t�S����dV.�i�k��M̭9�!�g4E���I4�t�����Q��9�il�&��<���&ı�������2#�L�E�*r��d���A��S���@��Zj�����89�� e��b/�=��7?�[�.NR�]o��$�T��o���E�?��[�L�]}�p�[j�[��	p!k��ӭ{`I�<��j�=(f�b� �\#�g7[�h����J������y7��Kٯ��_cE7��xKg!#�v��^���~�Ԟ���XX�fT�G*էX���ܶ�0�x0գp�:�&�ڠ�㠀b=28��
:�ܾ�K_S���ޡw^a�f��k`7zl�:���[�����b"՘�=e��z`��o��2����Tj�Z�|X����ߢ�AX,3;	t{��2�����+���lU�­6Da�؇�R�Sy'��=�]�%*�l#
�L?`v��ꞷ�G
+׫ln�q�0�����PPp`��i"+~�e/ʵ�}17*�Mײ�-�W�u#�l??^���4PO
t2!�F�+��n�	\���c'�bp�&5�������<���q�/��
P	�2Dd�'$~�I���ޭ�>�"d�F?�&
��Ӆ�H��D�
+"�5O�V��͈�x�9P��dh�)0�޵:�C���X�W5TIw�l�*�I��.�RM
�'%$�8��\�Q\S`��cG�jK�@b��P�d\{�Po�����USY+y���H���eS4�ά R���d3��>��O�l(g)U�h�Կ�[;ϛ�����-|����ΈŘ;oZ5��;���d̦���m�5Lul�׊b�ٔ�7���舘*��a�����k��>�W�ٴ|�K>��p)P��x�,�GG\= ��������U3 ��%ߟ���W2BB~����4���guXګ���1��#���L�wV��o�E��M��hBz����!l�dm$��8"��`c{���.+�?�M�g��fbv��B��ro�?2�8�SS�&Z)͎�D��4�h��tT�Ǥ���XY�a��Y�[������������K���d"�^&cS�J�N���1c=�4��YԚ"+�9|�ؐE3E���Zi��X9���R\��~w�R����Af��Q��H!�)(Aӟ���k�v����J��]��4o%@�����Ut�܂f9��=�+���hz�W���Mz�ǥ���X��
Ӹ X�t��m��f�����U���w]�L�oS,�#�$5�d7��#Ύ#��B�o��մH�m��5z�6��*f'@��+/��#�	Y�ۗ�I�w=�Ӛn7�Y�Ŵ*\�O��SL�c�>�Ulд(��%M�7��>�V�'?0�l*��ȼm��&�+��k��erL`���W)�x���Ȋ���M�-�%uF6t= !��!���n_����x+��G}M��}6��X�m����ٶ����5yٗ#��f�1NU�^d��Ƭ�H�E��a�ƊM�!E��E0ҁ8�=&϶mC��+&5��}���kp&�hg���^��Mh�%	�q�ڶm[I�ň�7��)sgv94{����e��6� c������y��S��W[D�/��GP�̽� ���+b��Өw�x\��>�= yba�|�/a�f�n3_\�:��l��z����XAt�t���Y�:�����|r���\�q\,�}+���In�t��J��Fy2���8��ן[��:���i�oϙ��j���X���n_;,U:�Z�Cn@��OMH���-Z_aP��-W���t&|����G�J��	iQH��6Fb��$�����f},�j�C\�*L�3��)�����iI��aV��3{�i�ALڃ������a�>5���v/����7���1�t���X{pɳKʠ�cÑ�.� ��Y�g���ka�t���IH�K\Mc� ��+d�8Jw'��UT���}/��J�qy�7�6�T����
k�-.�aP^�z�i���0����^�I �7�Cb��v`�e�T%�E�H�g
��h}c��W����Sr\^��o�m����P��L��ɠ¢n���ê����[�*㪒0(9o6��ª�v��Vb(a��=p�DBz���� b�f��!��.�R�/�(�v�P�4j��Ufy�]~��[�e�o<�5�v�̘��zu�J���\)���*���Æ=��I�%�t�d��8�D�a��f�#�O32��:�K��V������)5�e#�i��2烢��G�j�-j�)�j^��7t<6��a�V���:�p���5��9]���Xp��nn�m5��(��`�9��3OBrDk�Q�xؼ�n1U�0U�Y�Ǹ��������^��?ҋ.Z�V���=��-�B�QC�K�w���E�ҿd�J7r�0v4���[����`�h_ 3�p�P$�9�JC׳���Y�o����,��k�Q��~�Az�.c�-2tG[,�AE2@�%�� _ �;�n�Ǽ�@��g��79@�A�p��n�E��D}ɥ���w���=wbSk���jEP�3��Ϗ� ��/m�7�֤�gY'|��x2L0��"��нL����$��F)�]G$��E)��(���V͞�k��q�IFX�$G�j|��,9����(d�p��"ɷ?%�݌l\��6�}u��(w4sm�,�]��_}R�Ia�g��\�0C������a6�`)!G�Wx�P�ݗ�G=����Y�i�r/0p`�pT�Rӏ 6 �,��\��~^�=o���;��^��XN^��7F[���uU��3z\�P�kfI�J��B����yC�/`��/�d
%����Б���0����h���+}���8p]��P���ě��5�+e�?�$c�ET������<0��Ā��nh`�NǏ���B �;9��;뤙j]�.�+Ei�7\N��F��	�U�3@{i�ftg�^U�檈�,T�NE8��<,�i��^��V��\׫ԫ���;;�k/�کIF�I���>2 C�^n�)`��xCGeW�@��-�T�ʉF�l��Y����F�ER����� �}��YN�t�	�|zDfێBGl��52�v�s+iM�+⏘�����Y�}��û�����~�b
4[m�uƓa���R�j�r���@ŀX?`��P)g���l����n3�����(ʜ^�X�l
�^KS�Ϗ�MZ�y+�j�򽒓�.+��x�/�C��])�l���Z�4�L�To�v1��Tc��R  �iMG�?��s� X{�M�S��*�t�����t��v��ڌ���ϋ׋)k��;�UqY�S�q\1:VSw(O@6�`$�(��n܍�!��O�駋/���}KJ�Β��S6����֩,�6:ƈ:��g|�*�M;s�(ާkg��;��*x��s�Z4(IF�osU>'虖�����Dе�n�'�l�ɐ.b5�bDÜ����ke�`�������䁀�HމM%�h�Q#��ȶ����/�;�F�T�R�mM�h�$F!|��jG5�
�:�LIo$6�����J�����r,v�=��aGy#q��@$��N�]�M���x�m:�[���F��jw]�R��Mħ���y�-1A�v�viFqe�� 	��%N��JJ�G"���X��b<^��X�U��b�&��l���Z������:$F"���(�Z[�\��s��c,��`)=���"��͠�#]�#D2f��P[��cw:O�����)[�j.�n�L�*���=C�@Y���U� �r� H���J�u����L�1[������񉾂?ׯ���1rb�+DD	��9��L\�+�y������6�x/��`����`�E.]���R�,������$�������l�oW �*I��?d�p�6��|���k[WK�����K"%�U?�>Q;>���'o��������p�&�5J��K��tp��\�d�K�22����@R?�ܶ��tI�#O�A��h�\�G�"��R,�~�->$FmX�}���B�(u]�۶��j����p��qQ��~
�Wh�6�3�^�s��!|3vꤜ?�l��
�O����3q��w�J�l�C'��z��c�*��H�$�'z��S>P����{���[ ��R��!5C�&�"�����șB`B�E��S�d_Be��V�^��Xvv7b���/��.	�L^��(�+���˼����j#cOx,w��:6
dH�.p⬁�}�3T����q.\�J�7P��Rd�'CΒvq�j��K��/P���
]^6��l
i�&k���8��H�DI>� �Sb�����0|2@��_�������6�Z��ԋ�{t�d=҉�<ʷo�#�"cYh+���(��{$�X(�P+��N�a6��EE:��>�՟�) ���"u��ƚ�t���#�Ƛ�\��ׅV]K��<\렅��/�Bd�5И)�7t(��{�^\
<�����qn�����RU��e�� Z��1�O�Ve廖��(ح^�5Et�X��\9�4�8���g ��N��	��2ReY�5����K�3��Ѣ�y��3����8{XY�<�`�d٥����^���G��x?H�,ROA�!���-�D,�P%�!Y�-���ܰ��L�	��N�Q�fOkL���N�[�o� ڟ1��J��Phރō��,^& �V��x��E��/5x�����u���t���K!����xV�\gԸ:�B��DTFk�EX��nK�ۃ��>��X�J��P3��f9�����_�Ͷj�;�>9�J2ǷE��l���ϧjw���*�/�N�F����&&�>��YH\n��pB���t�$ ywf��+x$��{�n�(kA�de���rM���"�����*�j  w�_eG��'ـ�����ta�u
�������&��������LD��2>'���:S�s��l/�Mױ��,��;1K!��~5�aG<�E���vr٩� ��Au�;rC����F�ܫ&>[�	儳S{C����[1m��� G�8@�Z��IG�� �I��K%���+9��&��d���c�5d	�ߣ�����~�S��x�����t�"g�T�h�<I�C��;f�y����͈ey�MH��e���^��Δ9��MF�*��������ً��S�����M'
���{��u���c��`j9jb��Қ�XB,�����:b9wڍ� 1��Aaܜ�Ǧ���:�W���ML��>S|����9���T޲��Q��$0&��s��k�ґ>�7
�;��&ͅ�1��3R�ؐ���I��j�U��	R"���@RaJHO-z��L,>�[nƚ�>դj��(�j���h�=����𒀒�5$1�B
Bzh��Dۘb#]�<�
׸�$ԉ���}�H�\.��RV���V�{4�e�E� C�.!R�F}�3P���T����p׫D�������4Rr�f��CN 䮞�D�Wh��%Q'�Q��҃8� yctI��+ Ҭ�f��y�������HR�L�{��8��@�Q�¼�2SY���w�EcV1Q��t0�E����J+���3KXXZ�zx��n��h'�-K ��m�w�g6��>�z&��_������G/N����$$ �Ζ�,��j>a:�D�*�pu=K�U^����Վ�`�1����s�YP��S��,2SR�ҏ_tk�9,�iT߶
�<���u�j7b]EL[�Z��.XG�im4��9��X�k
���8xi���l8�u0�`��l���M�/GKi��H|:&��(HMսש�G�7��/�e]�������Ξ�Ʃx�p�X�B�P-�����5�B�Pw����p��� �ͯ�PI���>����>2%�f%��D��n�P�J��|�e!�4�Ͽ��3��$]�_N�(g*��0G�c��C<�3�yH��f��b��T�4:8&�pH�H�/R�جxK�X?U*r��n���]�瑧e�|�6�]��g`�COۖG��et/Cb��*��}���;���&!`+��V���	~��
������wj���ڏ5*�C��>������� d\���)��vS�H�[���;�r�4�	���7u��P�f<��U�2���ь1�%�11� Z&�j�1��Z����V$?��eD�2%�O�x���)�|_-	�ˀ�t+0�*K��)G���6�YX6�(39,�������q��b���u�Ϟ�g�4���]ʪ}�ĺ��pi���Y��s����@�4&����2aS9p����M��0 J�i����($>���
����8�d�"&4�����:h��!�&oK���>�=0�#d3@��(�� ����q)�f�Z"z� eF�ם�:��#y�� C;mO�m4
_͋-%}f�� 1Ll0��D��&`m��.,���+7+B�N�j�6�9}������gg�K��ܿ ���<��C�����^��50y+�	c�-��~�vC� �9� ���q�����6v�i�G'�@��O��x��E/���D"rw��JpV�{���g^��8�xg��A�*E"�G�ީ���3U�||G�S��&���$# ��.���s@ȋ:�K�;�RN��Y�a���B=�0{���%=��*V�F�nw8��HKd��@�,���# 6��������'H��i�������Q`w��0�,�O�Z��l��J'
�C:��6�](�k&\TҊ��iD9R:�e�����~04�ց)(V����1�oLX˴���D�����#-d�VI��ͻU���eK�*U��u���o��9p%�>R:�m�W�� O,�&l�n�����L����]���K �3��8��L�H<

ܐe�N�׍K�'��/���-X+v�;��,������+�k��6o�y�L�* �6�Q�}���:U�[�����U��s˦�46%&󟣛b�7�?�0{a���L\��P����>B/.�"�,vC���&�w�s�F�$������cݳ�Q,�L��)V��ܞ¾c8��E�љ!n�E���r�y�}O)��K^&Nm~��O�w�/�(� �]��\�f��iZF�t&A�	m�J��x��Uɛӡ��6^"q=$�O�Y������S�F*�lBd�sJ����~���X������f}��'��"`�̨im":E�N^�Z��v��o��Ky���J�f:�N�_yd����&�-Tۋ�ȅd�d�[4"����`}�|������v�L�"�eʹM��PY�;6�%�!�=�բɮ��x\���T!F65v��|����������G��Dc.�4z������-D�Y�y��Ni��p��/0�?ܙe�,�E��fNnG��\JY��D��R�||C�\�s��,����gA���f�Kx�]� w�_����*RK����⇊��L���3t
�O�D���=.F�E=g�\�l�m>�}ǌa���66@���ܗ�Ma�m�E��F<��6��TW�Ծ�k�0��=o\�ց�qq�]�Yϼ�{s�B����PZ���"0-#F0:k4ܬ1^���A�Ý��P��O'��8=���C��j���bT�Ŕ�v(�V���+��wO�5���D��'�$��4;�a����$���+�S��J-:�WϢ�V,"[�ԩ9㯶o�ޙ�s��t���s��v���'�8ب�]@�b��+:��o\:� ��v�Rh�g~�_Ҟ5p;�c\[%:��5eV��<�K;��liE�<l"�U1CO箨�X�{A�9��(�(x�-�c����*�h�2�⯫or~;)�Pp�Q�*ِ	�.�+Q/��ڝ��A�C�q_��Zd�^;���Nv�3h~��'u��m��?�}�k�i��ςbE�P�E%  d�AX�S�; g_m�fM�:ɲ��R�x�:9)�'.Ѭ6�a�;��D�
E�e�;D����-���]�;O���c����k��e�E�&��C�tƓ�$t2}24k�%���7l�ЗA�ͼr�.?��2�:
B�'/���?�U^��	��֜������-<�(���G�}o>$��"�f�ʈ�g�n#S`�e}wv��G�8/إ0Y�0;t.�y�k��Ta	�9�"To�,�{y3�q|�����jo���B�Gmr&���])Z�ڛx�g�[�r�n�b]�U�35}�h�-O�nH���5�պ��x�M�^��JVp�ky\��lP��OQ������j��03�t,��!-�q��My�	�����E�����y��/o�!�g��	�)w�?���k%&m��ֳ�������i�����(�`��_x��&B�L�*���FN�^��Yo�l������2�-�{�4���E؆��#����ݝY�_�Y|�6��?�nc�@�U��4s��~�q7<����H�*~�f���������緄Ζ���9���BdU\���`�M��R$]Ge3�c�@
6�5���#k����03o�XV�n�%�-�x��!��Q��.p���k#�՜2���f6�҃��4]�H�2p���R9�Y>���a����J<��E�V�h���2x�6R�Q)���kED��xҶd��)Ri[�~)y�	�ڏ��\��i��k����J�d�A^�;�z��4�p���bxh�R��S���-)8���{U�ǭ
*!���0Z6*��^���?�V'���� �4��2X='�w;�!B�eU@O�����c9�����kr�2�v!�9��i��h�����"�f���w9�,�H���xSjD��<�����v ._C�vS��+���aT�x�fe��^1��y��F[vx�{ѳ^۳G��'�O?�%:L��x�6��{�z(_|%�� �.���C������_���ԭ1���v�A��W���H_>�ʀ���5�������g�X�{f���=8�[�?L7x=m*	T�6�'!R�s/�c���<[�[�Y���j^��0ϭ��VY��!�q>�0�툋2�EE�׀�j�?������lu�� %��_��j�(��H �N`m��/s�C?ח� �f���u+C~�cȶ�(j�%��^�M+�c�lC��mq�`���7��=	���}�fn�o���BCt�=z3!�����j����������ᣂ������"b�3C�:���9�x+��9~S�^�"5\����Y���^+�� ?� *��[�T��3���8�D�l�f��i��d6�%?��.w��6���J���r|��]U����g� '�����;���V�+Vj��/X�wl�t����W�3~Ќ��/�}z텰XI��Mຠ��z��7O=���$G��c���ћ�yBbo#f�aV�Ο�k��6��\WНOC�RJ�p�q��G<{��p(�����`���;����_/%��}uQga\�}��M4�������/���MI�3d�ų[5��PV�hԛ����
�^h�!jǦ��yz��ߣ��V�)�s�?V��R<Rf�����%G�[�J��$t�{�Y�u����R,��.vA��*aV<�g$��� ����yf�h�ܕ1R�t�.���Cʽ;��%WUe����`���:����r���
d�$��B���*�f{ �"��jLviB�[V�	Ķ�u��P�cT�x{U�p�G��afi'2]�A�R,>|'B�!^�_�\� U���=/�Ҩ%�~��&�-�=���!�]��+�0��J������)��Yb�S�gX���R�,
�����4XH[[�]Z&e��q'yX6�rT�A��x�z�yz��"BUD�v|v����BG��o$N���;秾�O�n4�=CPԐ���E��r�W�Hi�DD��@~���.�)~
2ty �Z�n��'!,F�h�Ȇ<�������������_�긕�r!��A�*Ώ.���ދ�����O.�S�����o\��?,���������_�0�`8͖4�#=��T�a���>T�#�6�`��R�|�A����}�^�߷��(��|o�-6�W����?!�y��D<"��q/�����_�J��8D��؁�]�
�gE�&�PA4r���&�'q#��!������θ��hyr��Z]`�r)��L�҅]��2!Ρ�C���
6g�$/��p[��RZ`4���4���? �}�
vx�l�
%�>b���MW�9��a�zX�)�@�ˆ�c!��~��c�X��6�G�K�)�3ͯK�(3�x`|��o��䯯�-��?��'��W�/ ���@��ު�Ȳj�O����s	ܠ##��j�e� �d��77�I�p'��S�l�C(z"��p��~��2Ц��.`I�aC�9�vFl\l'�^�K����6q�e� I���}�h�@��C���YF��H�MV��.{�[֨�Q_?8���VGm�����D�f���Y�|�sՏq�;Y���D^�>Gط���/�i�3��|R��^�/mc��Fp3$6�a:ѡ�k5*���n���+q���Q��?ӯ�p���E�~v_��"G�E`���� ���m��#0jM2$��k/9F+>�"����;�d���k�Z�sLs{�L��y~z�Bլk�@�6��בv�4oh�;�f�o���OS�#8,n�����g4�i����5s{a%'~��T�	�~M�1 �黟��]�%�Dގ�����`4�}��d�I���q���ɮF-�3}��n�L+B�d&�ER&����r�f*�� [sJ�a��?��l��j]�����ڙ�h�����������iý�Τ�b*oc	�`�ӓl
%�O����_�C��v��slǣ9;{^԰�A?9����i�Am�#�@	�	`��k�Ƅ��csj�n�O3�S��ʅC��Ɖ����Eq_*�ha�{�9V�Isezv��z�<I9.`4�0��
��9�ES�ߐ|���?�[9ݑ��po	_xN��K��d��X�m�N�vԬ/���i5�5�ʿ�v�X�X���p��1 �����'g����³`���&g�@��L��8V�g���Ŵ�К���Q4�@�8�ZJ�$xo�A���_�ga����Ē�X��;t�5���4��ܧ�������3�|�z��	��%�� �Ҁ�r��4!�j�<����0�G|�-�n��ߧ;�nˌ���S�G%�0�y�xB��|1����&]�2/�R��Ѕ��՗����y�9���~�
گ�M�J����aε���P{�̈́2���c<��H]����gg�Ѕ���[3��P��&Q��2�;1B�䋹k���4�Aļr�E���I�3Rr}��.�	�d���T��1��i��K����:���Z�b�������>"�C1��1)��ƿ�KR��[g5��gT��
���~vaHތ�⽭��b�B�J�y�b�֥�=�<S��B�)��^s%m����$�_��&�ܫp����Yy�A����o�+�Dv�̣
j|X������n�g{8=���!!�sJ)M)��������$ӹ6�i����Į�7U4 _AGc�ֿ
�j[s��r�(��F�0����Y�^j����8��)(cy��z���[$z��3r�"9_�sdD�F��_�@,0�)�>␮�w�x8�E�6��G�] [8g����X�.��٦�KG�(������0UV|�����`�m
2D��vĮ;���_�� bJJ1�(c�/�f��q/�L..�"ҡ�e�>^�\����?���#���.T�}@��_�̆+��<�Q�X��G�nj���{V5�8�е�j˞	���׉�O�[����"ܙ ev��b�l��<�{�?ƨ�y��nc��n0��	�� (�X��L�b�1DZHU��1M�)��e��^'�u+c�1�ڇ,�1�4�ZlA*Z�EK�A��۵��8�ki NXcF�o	��0Ö�Z��I$T��)��ա֨��Rh��j��(�4��*�n7�/)eT�Q>~�0p������GY	j|;�̎w�+&��{��Q+��@"\|`�����G8,���a~���\��hQ�$��c�C�8�o����X��t;�j#�V|�ǃ�e�����[��Y�nSMZa2N���;��}�P]	���ڌl;bE�3BoNjQ�~��s�2��T��� g%�a R3s5M�x�MB��a��t�����I���b8�� i���hi�	u�����uA澱�-���-KU>r!��ȚB��S�55��kJ1f\V�-B����:�}��q���S������氒W�9��=�7f�,/Z����]?�aЈ����1W��5��o�F�a�Q㤶$[�Ϥ>�*��ʞ	R�Y���o�� >�����)�!�n��'=�U�t��ݬ�d�xB��Y��a�	�����)��TVޠ�*�xD��]I����N���z�'s���wpԂu:Q���N`Ӊ��9>Pw���<��A�ʚ9]c���1�TCV��R���(��cb>f��v4>tpS�N�*
9$5R���G*�#~OR��<U�;l(���Fr�C�bK�}m-۰���_MC���q�����h�/7�{*�[&s��i-x��`�B=��V���9L�'�ߎ�V&]�Q���ճ��BE�'h �3�7-�v�H����|{��*�E�	,ba�_��H�S��n�E.��#�V�[�f��y!�h�U�"�@�zt��/!�k�Ðj�F�B�
�)�
V�� /`��'S����p�%�3�>s�4���1�,��F�8��4�.4�,��w�,O`3,�����!�w�=^�n���aQ�)������g�
>�na�&��,�,�Avc��y�r�9���`o^����е�]��L�E�ĕ���+1������+�p��1�b���*!������x�e��x/�!�e���5,؄����������%+��J����nײ�Sy�=���]Y�9��ЁQ��G���?��cΩCT�9��;Q*Wl�	r2�g�L��\�`T���kW�G�sz<&��v^���1��V#�gyC� �h-r�-Oת�,z
\����3�yɜ���^(�T�F��������;��J-����)�#�!��+��?J6h�죺?�g��ID���`�4��ʼ�t�؉}:5�x>��<d����t`%�����(��;�	�����[[
�-<��q�. �"����Eӫ���c��ߤ�)m�>��F*�y���+5GlB�+q@��0쁺�D�WY
>W;��P�W�Io\� "�c!�J[�n��z(v�9�K�W�����+�e��9����\5wO��m^K�?�-��L|=1�4��T��I�� ��"�u�e�߰�h�J�?Y���Zx��vqf��7� y2nۯ>K��!���)dF�x
7��qX���b\�$Wtn�2.����c�Vțw�+u��#=FD�8-]y<�,�Ɂ �Bw����>ĝ�J3b��ˏ �W�x'��A,}L\�8U�r� ö�b�7ǧP�������^\�QO*;Ap��Q�r�ϵ�?��_���Rf*S���)T����&��X����Jz��vާ�@��a��0����
��@-q�	�b��j:���l��E��ޓy���HoL�-�0��Ǿ���mwI���:�<HI�5��Yl����q�	n����d��oY�GȿO){u����
��Z״~�`�Ͻ��ܚ'Tx�=�(��Re�2{��1�g롤�@<RH�ʓC�ȉT�G$�2��g��t�4QG��}Ρ����9v���D#h�K������9G<5���kMa oׁ�0ħ�eY��kgVYlﳉ.!�h�bkd▝ar�����h�2���aҦr�jA�@�+�����#�h/�w�'7�g|	Q7,��t�:ȌS�[��|��rǞ�Fegt��#���FX!7�D��3����B�c�M��-L0��Fk���W��P���U�`�l�<c�:R�ԼoH����R9<b���N�%ӈ�#����p�鯎�c��� ��d[�\��"��������z�M@��F��8?�,�7�G��p6aDi�y:��0i�a�P �l�H�����J��˓&D�a�]wR��b�	JVNH�_ �>�Z`\���j�k��������9�Xؾ��@
�a���N�B�".��4�6�N���)�i L8��\|8B+��C#j�4_���m쉯�$2ul%?[:q�t�N�W��9�?k��o�Ϻ [�`dmuސ�IQj�{�D�4oT�wf��v�x_�^�Pp$� �e���d�Уq	��ؕ��ą�Η�|"-�i���?ϟ�����y��+n�6c^
���%(~-sF�E�U�0�e�j|h����'Y��<D[��:ߧ�Ue�	b�s��FcpJ_�.?7X�A�P,�2K:�W*
k�����f�����q@=`�͈��o���Yx�,��Uի�i����Y�7H�"ь	rMϽ���az�Ǐ[#-�j{tA>ڰJwGk��˞��U��.���U�3MW������ iA;5��H�s"'٠���L���8���-����^��[�L�aˁk�@#�t��l��D�����^	����U��q6�L%H`=¬]�N��J!6�;l#���rΊ���(��z5k�t�Ӓ�¥�\�8���m�K[�ia]\�>y�������bWŕ�=�����Z����M�e���(Uy�>���i	����n���.�?������&�Y��I5;�������v�w�\a�˙n>��<U�TTRr�KnKW4r|��w�Vkp"ys��ε�@�wu'��!�C�@YcƱ��|��c#��K(�h)�M� ���������5���y!��F�i����nRٳ������p�/h�7wƱ�/���i��TK�U�n����
b�@qד�gP�$�H�Qi�HS6��bJl�
�^�<as��j�g� U��c������BBH��$p�m#,�R��bh��Hq�p�-bX	�^B��hNU8�&��L��,&?`��5��l.���� ̭�"�lK��g|�N�l�s=K�^s��0�gLy`�#��ֿn��Z)<9	�!���x� �뺯�{D�[�2�Wyƽ5x�5����e�K�=x��ް�����Լ�Zx��/����n��>�m�
�ҍA��g�Z���f�&��l��4�*Y������Q������^��ׅ��H �h��N)t�����cs�[f���D`��g�~�� ʐO�Lv���av�C�����z���}Q��F%�^c�J���u��_K�QD>�x���ݘC��ݏf娺(;���sk�S��5��0(~ �p�1��5V
0N�D�9��*9: 	���u��^S�F����x} Y劒�оjH����(�Ѧ���,�C=�-0�E���
��8�Ht��FT��Ĺ���'�-+����ɪ)�c�W�m��(����D����qA0�mM��]E�����f�*GP(�%c�}��c!���=�n`̻
��>�o�8��/%����@���J���u�q��O�����^��1Zm����1+�7�nd,	 c<⑨��6���jP��`i ���6��J©hv�6����0�y�I-&��ʉ�d8o�n�[y(~Ț.�Hyv3E_aP33�N�_��z���0L[�80��H�Z<��k�/��J=���h�� �$~��$f�Z��5�ĸ��*�M�LSs�]Z/��T���Ӫ������l��[̙�����7�#�K*��;r�W'�hW�X���8�@Y���3� =�(��c�.�&NخΆR�]<M��oŞ�pu�f,؉o���Nj\��q���'��gw2}�N,Ψ�hS4��T�t��,������ZSt!}��Xvyv�L*�B|o^@������bh���Z`9d�������~/�L������]���:��V(q�Ap�����ɪ~ƢbU����6-�R7�S�=/�������Q��ae�'�K�l�R�#!��nG��&DC-��4�*^��l g�A���E��9G�� �+�#��4`,�x���hD�=)�<:zVBZ��1j]��5@��%Ke51�ԧ�>ۚx�&�B;���z�Q:�P������{����-~�J� �ޔ���å�L������q1+�$J��(�~��f�l���m�Ru���k�1)�4�, s҅���+�Y��=������Ϧ-��\�IN�7�rm��-�>����@ziN"��!O�P���/����g�FԖL��4:��3nn�16"�o$�����^���V�F�P�+�X		�[`@��Q,|�^�>�TM"]�N��A^z���V{wo���]���[}I�&��f.�&�ؽ0���4ۊ*\`�ĕʱ?.��<Ť˺dzf6;x�Б�����P��+�?�>���Ɯ�}�K���Y�ʥ+6p(^V�4^Lr��&~��bb;�*Z�-��`�IL��gl����\��kz�U�d	ɟ �)�����oMo{j*�M��JW~��G�}�������hԹqqΉ"���&o���?ņa��5~U�'�!��i{����}������FS榫3�;˻k��Rh���1^5c�5T��[:�l�!)g�^r����;,D�=L��G<<�e;IJ(���_7���÷�. ޶�u&xm+�J��O��:�r7@j�X ;rϵH�¼HJ��@��*�!����bQ�2Y��W��>\eӉ_wcu�ߟ�x��].6�������`P	�3/��8Z&��^?�a�Yڠ5&ԫhp	ֻ�5���W���Wd}�ۤPE����rNfiͰb-T��a>�Ϡ])�?N�iv�P5�=!b�}�f4i��9n0��{�����-?��;lت��.�3�s��p�	����p� �%8sq9jW�3��J�O�׫���e�"zǊZ�cG��c�K��߽���6 �kc¯�J�pLmq��E�+w�����o�����a�[#^'Ln0q�w� �+,Է�ooO\��띹	���6���䥱���-��.⍰�[�0c�3P
�U&7':_M��T:����^KD�g�㶜b$K�b�� �4�q�!/
�g]�E�����2U����>3���)�T�������D��aa�P�\�d1��qx�NG�`�&����=F ���������~R�0'�*s�9�?��8��'5`ۛm������e���!#���xB���W>�����ce���w�V��&6�u��5��Lw�*]4��N,1��|��X��M¥n�h ,��.�|����:�gS��(3��!h:��y'-��+5��:��U?���]W�kP'��6��w�G+�<R_��+� $$2��z����8����D~�_Q���/D��Uqwk�F��sn5>����1�8�I�m�rL�]��y�6��N<��v��bK��I ޏ�����w
l����&����K`X�'j��vl:�͝р�|���B����	3R��{j��U�+�L��w�۩���ڶ;0icܱ�_��2Xʍ~t���;������ៈ����U:�!X���F�y��T��e5�|��nO纋Qɂ��b�x�-g�O���j�_n�\`�'�Q��@��͚�: ��oA��^�85�8�ø3v�h%������ȼ�5���X�I_��{�L�������I���'ϴ@)n�c�0��岶����*- �}:��vܔ`�$�|��?,�Qz7�{�߁�d�ɑ�2�v������K!!�*s�� �kd����nD������y|�}kƨw�B�-�i�R��7��˿�H���u�e#iW��3-�<�DK��}H@�Y@O�΢�;�hd�s�`��`� |;F�}�;p#�*�j�S����Jd��c�,y��p0��.)`G̰��F��HdN<tN^�)�\�;��@뗾��	��A��Յhʅ�~hJ�o����xht��x�I�09���*}(�L`i~E��?c;9�����+O�����`�x�Ԛ��Жn}�8��/!���RS�a�I'ov����	��"d^��X;n���_t�wܰ]�\S)�ʞm�ՠ�����퍾��io�Z����L�hװ��^�/��fD���v*�᝘ߧG�d���`�����"R�d8s���.�(�j/�@}���^:1�\��ds���O���x��C���p��}�O,�e��`^I����`�o�.�e���I
)��)�s\�H���*���M������gF�՛4�6r\p�d;a�<�sT# XD��h 0F3�]qJ�J���ħ�w��E6��A&�<W�B��p���֜b�B����vܵ�_p~s��E+;�/x�,�+�pؑ&G)���֔�x�V���<�S�"!���@i�4� �?�wT�jwyn8ؖFmƼ���8���Ƀj����m��1�ܝX+)��׹]����ӑ?P%������{�{!#-~�@�����M����yx��>��ȑdm�q:8�|z��1�(����<��Vd%�k�&�,s�I�b�(�^�Z����=��·6�W��p�Fi�����Ž�^W�T��_� S�S������qK��Ń�e��Z����䤳~#G�p1�D__��8|�&��l��zZf��3�"Qx�_X���Iz`\�AK��4a'��ϭ����@���
1�i�����jQ���[g~���,ef^%(����~"M���D,'�WK�*9����=��?��Dg&�_���<͍�����vA\y�+n���K�'������w�{#,�W��Ѯ����⠂`�#�3x�,j%�Ӣz��9^!_��m�9�B�+�����ӿے��!�N��Y}�����E·�zm:��h��8�=�}Q���Ӧ��'�w����Y�7P�3H�|`f-��Qf@��f���5���si��5�h>�mx�PH?$lh��w0�i�6�[�%�>����i�=�B�zSl�/�ĐTE{K�%>4�A�|�`a��9����#�2�ݿ��Fvn��"t��.N�jP*[Ņ"���ֻ�.��XQ���*(v@�.������˜�l@Ɓ�CW$u��丞�-��C��f���<�{C��D���v��҆;��X&�<%NmQ���-4G����g>�uA��hR��rn[�W����p��ŏ<O�p 7��zT֝��\p-0���{���)$]^��'g���O�,{3e;in&_`}�w�:��ZƏ�ڴ�G����!2�E�jv��V��j���5
�wL�;B~Ж�;��<y���z��7U��F�Ԧ���LM����G���F�g�g��[�-��:�"1����')���c��d��\Y�I��u,O��Vl{�xD��X�e�����P��R�����$���^rj��ޞ>>�yPΝ���'�hd?�I���F�e���n������M�#�(>�+[_H�^�4W��ed�q1�bmp� �,{�0�u�nRoK�C�R5��7������/�u.`�<b����L+2���^XI��b0.�F�ֹ
4�S�Mb��R� ;����יZ熾�1��z)��\���X�K���h;u��G�?�4\���?Q�h�t��,�����.�cbc͒�!����/���T�_�K+�	(��9�ɬ!�oP�JS�S��2��;�w��T�RUŻm�
[�Ό�z��3D�଀��S<*NI�\�{8�$g����J�m[0.ޭ����G�L'���#I�cI�ER#��˔c�o��"9�EhE�p��f���L�7N�4핮�!� ���U^�&�d[�\�����Itl��))���R}[��? +�dKa�n2H�<5E�Fp��т80|��)c�Ք�QDc����2�Ճ<S�aR����^Tu�jt)M|m��{r����U�[�����-9ds ́��3��N
'V��^P�Ԁ^�yG�{��T~?�Ӑi���(Jse�C����;��i��;��P�~�-�q^_�!���2]*0y���n�`B����lG3�gv�2b�plݲ�L��B)�����s��`��m�4�"%�a�`ϫ)=N@�4ieF���0_����}7�R�6t�E�K]� �j�X��!q)��~?�����ҒP�G��-��~�τod�g��x�y12�e��s�9�d�dC�f�I�L)����W�Chܘ���C-�aG�P��j��Db��Z�<�����X��br��xG��vd��Rݸ�\�������³Y⌮ʚ	��C��XBd���Z6�!���D	rw�h& ��+���'���'��d���Ѽk����hغ(f�����'��m/vӹ�8�nE�L�\��qC�Π����Xw����:Y:x�z��Fr�*����^xhd���ry�{U�^�;����R�C��Q��jt�����&��r>�Jl@iѵ^6��,1��K���	��������<r��J�y��9r0�������1"�/I�S��D��J�X��M��ĎE
�O@�x)����b�0u��z���*ļ�ᕡ�� 7P�I�*@��F��$��Y�J��5 �n�Q�*f�@y��G���Bw�gp�&]٨&RU�q�fL����C�q���V&Q������7`֐��i�ߥ}���ц��_-��E���&)S�P�� �?�����uaU�c��R5����T����o;|}o�M������!��'��!�Y���u��	v�~�{ ޔMӓK��ƶ
Z�ǌ�XS�+IV��"O�o�� Z7��7h'�
�j�w^�4�<2���h��ҧ�J�W�/��h9Y>t�8���Ȋ*�Q&�8��:8
�k�STJ1�v\�����^�"3~��6��쒺��O��"b�k"�O�w��A�4�4E�7�o������Փ������j�9� Hmm���F�)��g2�nxz�Q~:�l�Rs�����{G�����`'.u��툵�e
-�LjKm����n�M �x��[�[��f��8K�����g6�育b9v:k��"{�J����z��=v����8`i3�&Qٯp��C7�˙�SD�<^B�f�h��P�8���^�t�A�S���/U��e���!��;F�v��սwx�qx ����@�Ӓ1��e
�sS��f�c��Y#Ժ0��s��ϣ��g��+��(Fߙ�J돓��1�FL%G��A��CV��q��.aELh�/=�f���j?���97�l�m�k�}��G��o�ϗvb���bm��m[	��dE��ד��jr�@ډN��W&h��Y�j:���P)fi�N�A��z�T��ȡ$X��|�8b�	�D(70�x��/\���E#�$N\��� r��T����㯵�x����A#=A�Fn�d�v̟�Iz�|�좀�ej�axNl���w瀡OG|Q�-HJ����>�Hc,n�(a*���$��\�p���"�7��`�V���8���:��O�v�י���e{(�i�5����wjA �#�M��}ׁ�!�X�t�q��!4�{G�j�lM��S�������*���}D�C۾��)��UZ��(Jmu��e�jW��IbG��$�բbm�u����X�R<�ON
xR9]�O�!U � �=�-����nEL�Vu���;sD�=U��'qE_8�τ�����r��Ll�Au���Au��[j�M�ؙ3�7GS{�ӝ@���*�Ԋ���
��u�0	���ȵa~�>���'~3P4p�rgSe
�xWB�.{B�T��k��	�\Bjڇ>_OY�m�}�R�gb�b���~g��n8��9��	�I��-" �u1��HH���̓|RՂ�D΋QF|��N���U��h�Ǧ����Cޟ޿�2ˍ�M>V�Rg�K�i�2��Jס �֓%�[���R01ٲ�]bL�J���t�VJ�'����Q=n-���\k��.Q���]q�T����ӵt�IF�"��&Ԡ�".e�P)0��'b�zj/���y$��*���u-����`l�b/�mx+�<��PP���C���L"g�Ore���v,q�S�}�UZ0o���i<R��
q"�nQ���K=یp��߆���O?����	�|9�V�/�PIr?Lc��Ed+|�X�iF2�����c����\�������l9j4�4Nysy�%�p۩z����A��]�y����W�{�ᡐ=-�1�3�/���ȱ��()�A��0�ۚ5Jh��V������5n�go��8��9�H��i�m�
�B��.����\��`��h%�ٳ�nۘ�
��ш�ޥ?��ͬ[�M/H{��Z�z?}�k���Nu��r�"xD����<9A��1��D<��v������yU����>+%���2Q�uF��g�N��e6k�]Yh�"M�tF����S��/,�G�ɺA*pt�KX��Y��؊V��U�[$ ��"����[N��I�g�Z��M��1h|%��=V�\�� ��u��z�� z=�9#dJˇ��#��l�?w����YH?��gv��d�9I��Т*�!��+"���ŰƩ��-^�-���29:s���F�	��8����T����G����xqD�9��b�n)|�/%%��m|\�1��`���h�G�&;+�:��-{��5y���i��X�욨Җ�7�2|�5T�d� pb���+�[eow�Q���."'���W�QÌu�R�B��#��UKz��o=�S�N:���ƠR�����7����O����*�_±�'Ba�)3�j�ג��&�|��"g�Sq�ܳY8�O�jvoN���h1�Y*����� ��*����w�,���H_��B�a�s�qF��~�bt�&�(|a�z#y{)��|���2��Srg(�THԊ��f��/� ��Mdmqc^d��O���P�!�=�kvX�r]�/N`r���X\XH�%:��7���K�vy�R:���yַ��<dS)��_���_��Aڼ���ny+�7�{����e�tg�!�?UFU���۰S�>�ڿ���_���Y�r,�.pi����Sݥ�NYN�m��]�O)A�mq;ߥ��$�_m�S�s���Ko����,j��x_O�Rս��y��['m�x&�x]�y4@���Y[4��`Kr&R�ȱ7��5 �K��w�W��~x���ǹj 3T�Z��O�<��NrȨ@����0�1*�������!>cb㬶S %�Q�E�QA���2�ד����W�Á��4>��f��r���B�ȕ(.[(pg���sP�>e��X��,�=�ܥ9�IR����=��c�z�{�
K���$�\_�)Wq��R���.Nc�6�R~+o�K����N���.nÐ�K�r��+Aշ= @B��FS w%�ԥOK ��Xv+���Y-1��tG�?�k�9D���v�v�Tа7e�p����?tͺ
�>?(��#�����yj����޾�G�L�e��7^j���>�����5z��������#O�(C���7�Jn�v���|�߻�e�5x�/oE�9��B��8��
x�$U_{a�j�AL��}R���t�U%|����eb,��2�~Ɲ��(�(9̚����He�o�����JSf4�9�0���g�ٓU�zm����렇jG����F\�f���d�dz@��\X���>�EU'�
�3�p��5c���9~�O��7��1���(�j�Ȍւ��ͮ����"�er|bb���%2��l��,�gV��ˠ����mXri��k� {�E�U	��Ű;B|�	JP��o�t��_����D�T�"�� ��|#t���8�S�|�#�����{��o�*OXokt��������7gOoy���ń\�>W��z����6�qOE>J��7[�Ɔ"�2�Y[�����]��8�$�-OP��^E&͸L��+T���N�jp����ܽ\��x���#�3�ÈV�g���p>Yo.���*�;pD�ϼ�d�֨H>�����y:s�Z�h��i�0Svh�GwH@ʺ�q3�!c���-@; ��B�	M
��н�3�����j��ֳ�٠� 	����"���i2�O�%߶uȤ����z�����o��zJ�,X䟁�	(�P]B���nz����r}+x!�q�'�eTmj�I�ٹ�<]�3������ֹ�Y@wY�}!p���G��z�]!��ғ��׆T1>�{�u���|ͣ��F4�rM�Om�F2���_R�D8e+���c�+�uCYp��Ö֒�JE�G�,��B�ŘM��N� d�%rkU��_���2h|:��%iK�aC�.!f���h�ClGN��-���u�l�k�EWI��y2s��Jzvv-��һ��K�W�X�]��9��e��4�թ��\	�ܯ{h$Rª����(�\"�)��K�tL�V>���4�jHv���l�Tl�H4�p������]�T�;�{Pk��h���.[T��c��旙�[�RN
�����cLٳj��R�X~�&��Rs�u\��TR �Ύ>��i �s�z\������
��{k"<}��9�b�:�J�KT�+}H�W�� @�k��9�6�?�9�����v�C׎?�QgƒHv6e
��z�D��VyW�p���;����'.pn�-=f���IL>�|kE>����F/`g���u�`Ϟ�3_[�T�p��L��cQ�#�����I�B�ve)�ݎ©�5�7��yY�T�� ҦG3��
{Z惬q,��?�^1*D-8V�]�9 ����B-��kBU����Y�:=z�7����+��O��(���_r����~7���:����> �\�ڛ92e���2� ,��%;3e��#��d�Y�Aqq�����AϠs�`��������?� ,]M+�:�7��0��������T�+�����׆H!�o0{��G��x�zd��4���g}'����V^�J>�8�h.p������B���#|{�c��Q
�al�V\��?�*t銀B�r0����w�g���c*njI�O�Gs�j+7��B��@{��ݝ��h�w&X�Ѳ�xD����^>�T]蛈51;2Zb]�%��>�3�cFp�QF6�"��'�r��sy�n=m[����B���+�X��9I��޽8�O;PtN�z���E���Mz�&�Ho�f�0�h����Kj��"rs�n6�/|u�E�&\�j#Y9]��..����i��y�8����Z��mwNZM��Yջ��܇y'�v�~П�!��`�������Cdw�h���J�:�H������+��#�a�Tw�U����\��bEbib�|�8�@�o�
2!Żb* Filp8{gN.o �����o�s�������)�׃���V@��]qD(\̔�__�~�E{���Ȗ�����B)x�2�r�s:�D��0��k�B��a�宬]eٱO�ԚT���(�!��`c�2�0�����ۼ��o����$�����v;7�X�[>V 1����눚�!&J���b��:����B�P���]DPϦ\�{o�P')�T���;&K��s$������D0��������/��T|�z�:ԅ��9i�.pz* س�� jɍ��Q������:{�5:a����{��Qj�15��t���E k�^\z�&	~���p����=R�wJ�(<�(��S �]��&� 6����oXY�G!	���θ_���^K96�pY�iˇ��=2ڠ�o�Qݎ̈́�Vy24�����^g�~�r¦-��������m�iH�L�aL�{�!�əçS��*M��*ؗ	�G���6.1�x�~&�摬�ۑ���(F�C�C��r�� �EI���P�fܲ�6���Iܜ��{�UrƳe�kU~��5��|��R8l�Ϩ�5��]�����zQ��Lj��l�GIpئ��ci�zS�T�	�^�W�[b��Y"�\��d��e���E`�4���We�4�+!> /�)��|�I��]��P0`��+��DX��ѐ�L` cn�W�lʩZ(��]���Eٖ���|����r?L��%u��|��aP�[mH���V���m`BdNA��F&a�t,��oU�����a?u Ho�ed��e;�js�1#+�ʛ���p	o������,R
�*�˅��"���s��F4���WM�r�ϳfc@��1Q��id�LW2H�+�X���!<���H���zVB?�e��{��a�ÞN�z���	�/:�N:DE�c9���������.�*�]gK�\3��Pr8��Vw_􀌿s�Z;d�����-���,F�K-M����%lsD4�lUL�2����W%��g�^�z<�(L顛���ʲںy w?F#��?A���4�7a}%:���1B�$�Fw�um_������_�X��L�N���Fs#�[9d�Ie)A�R�?3���#n��[p'B�O�k}�`��_�>�輿�ߪ:���_<x:�=�P���D����f+�d_g~��Ի�d�⥵��<�ц�n�}t��Uڞ�n"W@�<�xvt"VHVȂx(K�C�L���F��@�8m&�ÊkTSw�����*G�͔�X�`fK<h��{٤�|�ȓ���A�T��曮f޳� �M[bZQ��C�c��l����f�>>"��m�"1�$l�B_��������,�� ���>Vsf�޲%+�e7Ї��'�UP,��鹥��s���w��#"Sq'u�iF�R�h� ����R���҉���x=�d#�j���^�d��sc�
������VXO��9sR2hp��b&tt�)�y���蹐�w'��m 8u���Y2?�,���D���ZN�EFp��)1��$`��p5��d��b̀5Ů/�8ܯ[�H�S�r��p��Ѐ���:fe�`�&����!�Qi>:U��i�;�� �+6���w�i!O~�@1��椬��g�Q�_5��JV][!�χy* >6����뀲L!��wE,薨�X�^|T��,�����	����ǿ��~n�U�w�֔SL�����3���
��QYh���1�΋��^{[(�jO �ْ�՜�wf��V�9���/j���m��{͓�wG[��,g��2�TnH&� �������s�� (��녕w��:�L𭩧C��|���<8��.1y��YQ���D��(\Wx@^�A3���7���+��tK���� ��3x
�17t��e�%$�کܣ�O~V�#P��W�3��o������a����$���k?�2��v�����%K�ka�O���#�W.� %k��?��՝�x�:+�&����8��U�P���"@S(rrQ�/z!��~� �_V�;;�Gv���Sӄ?;�x�İ9B�TΧ-���p���ب�A�).����b���y���	| ��q[�޾3T�C窯�#輛�Wk����!h�-Z^Wi���v���.>���Ѐ���Or��#�J�a�IOǕS1�;�çO�HJ��Y