-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
TLZojE5cdA20xvriQU80S3YYrsfVJBqox1LWsCaqfP0KyNMBA+FTWhYj8TnnmVNQQrnKu01H87ic
MpgSyqwAWY7baZ16RNRgEBR1SVNTnwdQmDrL38WSCzBu9j8Y/ktIgH6C7CR0HL4aCXmnKNCMv2tE
FqXTVa/0GEU/cv4+Fn+O6efIVKXCUFFYRHhxosnzSJ57hpIa0mpIoOU+DNOqx2a7yX3dB+5hbuLw
KmHnO/2WwOgPZFvbqMwCdgDqKbHN/avA08oHHa7qreI6NNBupX+koFAMP0lei/Wck4LKqdYbbffq
iJAuodMm5PbN2OPlXPQgrbH8FP/sQDEnogI08g==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 9712)
`protect data_block
M2722RI7PoWCuC/nOe9nDc3ZCCru/Q3ytVp0fSEIna3YAr5+iB9dyjIXdQKfp6h5xgBTUlYI/QVZ
hHkI6QKQ1wjYB/6XHZqCjY/AduKQW4kPigP3MzdHOKZSx9/6xAs0NuW2Z/wYZVtdOf6iieA7O2Yn
5h0nyzfphdOpYNIVpTKO9LUOylSnPKp57QkW2UCzPqFF3tqqcbpbENe5cZ1qsnQJicL5CO0dkvcT
laZTPZymroNZ5WKH3BjwidsOwZ9+U32zAlRng6/kTXhGf9djEUQf14+V6trBbF5DUxZ4arU8P76N
2uO1FZ6pCqbItcZfcV5B+h7A0ZYIHtikOTj06Lzy6gITTvC7cIUG8ERIZ3fgnpPN5ys/MwO75kGB
clqSobCemAq9+TaQjljEcme3KAKvPwtVIF0FQKM5MbqNGXapTd5YXLfzGJ85GoUvQeOuvOKFTf5M
hzV7k8HirwzB8eBWcD0KZg3ENwRxPvIcF0ea33hOz+BdRHU3+xIwQqsYLIX6ck7UT1unx5XX+kEm
Mp7G17IzG4iEN7V43P5GkQhlRxQwJoKQGPnKhjDXaidj2yz6MTsx7p1jxopvdi3Z+UP7JQajFsbJ
+pQklYT98w0/YuC0ThXEmFLqrvb+jOLDkjEhqTJWzkoH/cH+DQfPG5Sic4Qd7iWRn0Vvm7ykTBl5
oyB7Au9nS6Xc3M9K0LM4bRRSuG3PnWa3bB/CW4I9j8zCOMTODAQrxgh1Uv9A0qC3yVr/ZQRyIuyp
bPqkhndUv/jnFzOrYR1viO9DqLxhV28ELE6JStGvan/U9XT8DhvC8Y/gFJxNysiK5ZhM9d/r+fhy
4sziqLblNg7/5cEGxbU0oFCu3Lp0QXZfc531GU8bmfVo780aToMi60rTc0GZeB4N6HVL1LeeQff7
ssrfoh7o6nQ6yp78I/6srfG0G2MpNh1TMGJXgYgnx3YHlgttBQtTFaiJrz2AGvGq5/zWJOAypkLT
m7dd/TNuokrYipGvVcRjyhhfFhFOrcyGP3F9wWOYzngxGQNySLPy6WGqPqqHRl16xQiCDIcjfRaS
7JiME/FPlzEvt3MD6FCE1SdcUjJkSSCo4humDJqT/RKppmqADOA/B3R++KSjqO39Gd5mMgeL6Ev2
ICMmulqdV+qrLmKre69SE26xQhkNNULlxYg9qn5YeoFCxHAjJCF27Ftrkk5dA/BfenpAReqLy8eH
DAnh+r2NY5cvbByFWzfqqwDN095YnMJg5d4KZXzpiW8THC+82s+uqF5L2oVNxNTInk4BwDFYuYWq
N0JiIS3siuJpxOU4kn/CFot9g6vbJO31g/6+zuwI82B+159bwIvSfpDseTSga7sYbP/8T9i8B9cw
Pts0vNpeNoa3NF03iPd5tI44Gvfcrm2WHFbcTIdKc5jv4yqqrYtdxcZeQniGR+pvKGPtuTgpfN99
bP5Cs9epGpAyhCigTToJQmAShZwy48VywxojUhMlkZJOs4mRxMtVWL5irxbK3SrUzpZoF1vGbjqV
6INCXRYcrpLFSCiPchlcE4iWqABegv/EzufETNZWOrPj4nZtdTPB6L3YAipEvsb7F7ODcrKCWbDg
ZdtYo46/FZGXto1h/LDW65Srm3ai2PdgabAZ6MNfx+Gom4pu37bQrt1w6+06Lwd/Ft7M4ljQ0ZKI
Zq5nknPZcA5b9hTgZrgIOf2UDLjFv6Lo0JxML6j63R7QL1bj55GOl6NYIp6dKMJJSOvTj/ccNcq+
wLODM2EdvAKLagdRCYLP6uWJiUYa2CZ49U03nP5F96rbem84bTsdtGJgoqeIxRAac+oCC6evGv7e
8G9Pw4lp6ct8Jzpb4+MRVIhOuVimjFWLx4SQqWlRaOtF6HOH6G1x2JSJzsY0MIm70U055E5rSnJR
9j/u3ES8lTKpCRP3V5Xgj3PNSQDryQwWOZLE4ANHVeUWKZhc5zMH3LKQt8Z1/oEsM2ag68sYUCja
QUI7MJJQWY7WWmO14XuoJruf5Bx6YhfDsO93l+8zOmsrThuyl9mOaJOrDCxl18siBRy8SpRH8PQP
Lsgqxy3vXH+NU7p+JHh2jxUTtXnbLuXeDDfsGB+pa0AsYP4OxX8wn7G0fMVRqbgV3OtDzVa7nnCI
vl/qA/KMGrTeBIdI35GWkUddORwAORQ/z/6PGeOSzIASLRJ70V9aXPpJxD5f9q5PNji6vvqmR3Gq
KgQHo9pxKP6SERZmyZrRpv2i0RYmn2q8X8xXJGX9uIBAyMEpi7JqctEYAp4dfN3KY96RjQHiR3we
Hj5nnoNLexynP9VlKHDwBMyjEPvHn0dlcQ11GPnapsr15iq+TsLOd99LDssCMF69/JAVdfi5Fspw
NjQtzpWJtgWFqToon381wsrDxgEeTxVuTQ0vdQx73gzdiuBuf/GBBbH+N9A1sGvPKRm8kSQ7ptdK
i0cBZbWTZO+rQvIXn/XYnd6ufLiNZ8FEIAKqNhyar2bQGt5fXCI/ID5ZsDUAk8jYgI2mtqvUlBeS
LUXg0+F6IGUvHRsXty9Qf2iEVTK4GCTrfvkUkBcvOIRk8d6ugAAOmHd7CedcNQ9xg27kUqXs1YGj
bbRhq71XP7tceovHOGWyDydjJ6Pb6+gkFA8Xk1Y0nPKWzYsCR+xmFNmoe9VEmx26GMVQkBJUp38w
wqX/MGnc5AwMuAffuQ0fcz1Fs8MCQ1bwE8KCAt5Gc9c19HCrolEOh2OJLSLE03jxhAcCTIg/J550
rKUoaB5x3JMEQeMPlBdKQ9ypO+PXbzIJ/PCc64OTXUYwz9SyhWQlXSW+2SIoLf0cXpz2qQfQJLXK
T7IW4NaYYEVGrr7VVxWCQb0cGTEHk+7oMw1jnB6rpgi3VUPfJKB+2IwGaSb/hdwDdQJGkMAfutUM
7m2+j5nIiJrfKpXHIK11US0Kwd7u8ejcqpiQLz6vk14pao0pD36Y0IKpU7FP4SfWMth9m/bYx+NP
DVqVZ5A+kIkwo1fQc2QD8piJCXn+pYZ0nWPRctClskZxxXAMAQjT2Xz7ifVFPBaVy9NyMmTtAvRS
XI/H46ylGod1cOpWV18BfyYLij/2wDeoNRAXi1u48YWNicyi6oFJp12VdJzba0w/lzM+O9kBrV+x
lCm/Jq1wSxH9mpsnI6HVRUHb1gD5YWflaRPrIz1fQXrDE3yTb0Mlo1T5NZnYbzMhygH4ZP+vjL+n
6gVTiBeS5Fh91KDI88kho2XTRUqKPfmEy59HHKsbOSg2TZRVniiRekNYb93mD5eGMusGs1Dodesp
2AmS+Jraj6MANN5mdwD9qcwmo6yT5brAZWbnGtFwa6K5WwbCxbWmwWbcPsmxHZr1SzbazllBnprt
lm/hCeRgDnzKxqpFg2lZ6WehYENGvF8+0bERb/1dyUPRqGYdBKfbGBs595d50s7NeflQmFjexA5k
+4mdlMZO1VTXcqKROjqW/1+DgKMiQKMMsOEVYh8TZ//LRfZLs7Ayqc4AOpd7VUePdaMCdN/j6D8T
eYvyWJnNXm98sAiFbN/KRyj+ezBeYZnR0OjVdY8OmzKVbXq5ZnIEhRGcI+OcqvUBdjs4bFT9SnRx
5LRjnouFMAcE411OAm/Yirf05zBZHWZV3fvTrlteKDu9TNzL1uO5JruCvwp/Zb3gAJETROSY5tVI
9764Q1PYLI04+uc0vjQcguWNi66E3nOFEAgKByBrRFPXIwRzhBc3qC4wC2aZMinOdmydsoE+qRHn
fM9Z3jdLvYDC2AMQMe6Rpi8qOKVAEHMlwjyuwjmc65t+4lCm+Bbj1u4UikMI0gykXOhLWkHinvcL
bf6oecnBlww4znXp+GSxxceVd4qsEVVzCNKuHK7MIjR7FDiHFlhG/WnMrOFQQk7T1ZXy/WVhF3YN
e6L92+KsBXz1CcEcUKci03g6gqD3mRCnOZ6CTHYEd2k47skpuOwm8lKasgwl4baiWg+j/SdniciK
21XmNiCeO1M7KkySNiFyEAhbWtpPW4YkkiwRbnA+SaaRrortKjKcC6VsoqDToLiwmRrJRHPdIhtv
alBP0TU6MaH9Bhe+67PZT9VDb815I1vyMD1hYNeYcwYtZFvaioOwiRKInamVewhhg8fS6dyQtJBF
7PfjxdvCo4Fr6tUwUOPNZWvWx4+LtC/z/xX6AGtM61mpsXKEgjl3RTmqJuqzPHQR5ZeIDMXYaII2
a+G1exiwY3SLMgrjJ0aWjrTI2LMAArJqnhDvbX8Wb01XQsGBgxPFgr9coTUHFC9KW29A2akE3nnA
Od4tqyO8FonJyEUoi0ODxsqODWjwz1shUX4gj1Ough99Ju4Q8WKr7BZdiyvL3EDuaLVGt91OryGa
Pzlg7Hky4EE7yBEkM4QF8N4WVpetrZXnxNDBgwj4/hWvni0lEf+LbtSOFczNVoBWWC3J3tFBDzzM
ledUFW3S41ltJWQGQ36PKo6DV2ThDGXTTHL11J10L2UUs3z1CoQZyBHC7ltN4+fGaZh2Rs6fituy
QiKitd7VJRgkshgeq9ov4wvQcB6sWkGtv2rvpEqf3uzcCMiFi6NJ2jO69+mqwu5b5lbZ5kp404rc
72bKMKnCeM2QgTaHVyu4gYx1CmyKUbcNJEKOgFLcP4OM1lRuwhp9FuZGjpkFGys/jYX8pm6JCukL
t1vnH+zsArmtErvN5gxh2ueEIZmwaNTpl7KAEbyhLttNDm9wFf8t9vSM4YcB1ClORMj6TokARXdT
MePFopB0U7D7VS9AB2R90sPGX4OnYrf4BErjk45+enpvUSHq6H+08UrqBRaaNfKwbqWajJKIjTRF
Kg/iTVfll8bLz4eOqXrLvWa62/EN80E/FAlV5Ip5sC4cbDCURny8/xlWI57xkqJiWTudkG8ms2ao
M0Yu2Vp1Jhy4io+cWRgOSiuvU9J7SU7QSUay4FJLrLaGLKUgLLG343gzBsTD1y5eXJbGYakvalt4
yYvuskClBib01xOeG2e+Y7spwg/6MIOJQpYv877EM8iuaJm3Td5J3WjERaPUU8p2cWOSQsNElWyK
s7B/tBiLBxSvxFb297+Lm8z7nXlT+lDPhyHHwgP66PYZudEbKtSI3xI0YaJzXO8tA2OU3TgicT+X
dh0xPLe92Hk9CItRc6h1nhdYPJuBVydM7H+g0zE6LEUpHAmcZ61geLdvLGoh2NjtMc+qUdKi3bkt
zepzq29rY4+ZsNdfLhq96e4ArQaweQSoR58BcLujuUu29toDmhS6RovRWFrBL1fVsDiyGLqxlwOS
gO/fUHcTK8HfBtvcZiQ5QubfTH2Yhu5mZU9J5Be70zmQSVpDUXWzL2UD3Bz/I0EvcFcoUYnEQif2
y1xY1SK2BEjfhzqYOERV3IUr/X173uw2uXBbZUkCVlumPnXajGT7mlw7/RjvJ9Z7Ptq6xe2rSefM
KGnyKbUG9oEpYlaiELxDgILo8GjZ2oxug3H+y3GERpT5iPIeXpbTege9O5PF6FgzbhTMht7orG9L
OJUsSiK62bHuMo2aKmuh+oe3OZkRghcfseqnE05wrDM/xQkQBbowSSAmFF7sYf29T/RdLU2QgEHF
q0WAKywRgN/1vDc+w8T7rfyQjRazSUtlhQTV9avno5aJJLo6opO9mnjhag0fB3afk3dhnRa+YZle
iQxqtKarzANRYAqe+Yha+kS0evtmGvyiPLmKaYBapm1gODEjvGGs5SvTuTm+pBQ5qxOkbp7WPwHO
MnjbpMrDzhF1tfHmnnp19Gi/XE/0QRy40pSw5yTtiWSuxr5yWrONbeavyUamwWGwtyxDglJHvKDw
wg4FyOfCHZnAffRJS0M93XDchMumPW7iJm3y372+DsSRm/aP6fkLrbB9Em4TgJkDza1xOQrdcSfk
lyK/wm1EPTUe+uJI8iJP5q4x24BC0Jrthn5sXwypVHwFsI7fN9h2Rev36LO8wMkbWNRXAUKiLDy+
ncQl6KvovHP6sltx8qXsWdEJZwJ0SV7SFjo1Z8csdP0bXplqnLcjCJus1UqzwgmokyvYulj1X77s
Mt3bm3mi8sDVDLeoJEf53hrCPJF8Ag98rPTKHxa3I/QHsVwcR4z35SUz1i4L8Ppq1c7qdommH07D
Fzz6in6sRJD3p/6ecvy9CgPuoq+WRClwHP868lr+sAjsduNZLY8Qaekzn1s+N8sz0j/29l6BYN70
AOISn61s+LjjOu9sW2hpjRgQqgLxRMeElJ8uUQnDL1UFqdEItyEOSFYxlJ+eYX+gL/wGHK8Kat5n
m/LRhSjaEy6K4D1Lqnri5KrtFydEqpWxpGRiRTBXnEyQXd7yczoUZikJWb9CK6p3aYaQkaEOjxva
6lIsAyH2wgYPVOJ1x9VVG7OEoqHaFYoX32/46LmunKz108wvkAcsoKwSNEmtLna61DrVOobxc5Z3
0tNDXg4GKfK9PjY79aTIpNcbF/7aym12Rtsb28hS/A18B38/zCjKOADhHqUQVguii5wrAsg3NBJD
j09t9vWuMpo8BUPV4UH1g7IrfIRwsSKR3u57soA5G1Z8u/om0bNoF0kT6GOzsUadStdKcXz0p+S7
PzCjHnHe2I/CpHb4T7mpS0O2b2owOea+Sss28ZkqGU6Han+Oe9xDu8J2ZCxh8VQmrRRmAFcbwnLj
stFYftfRICs3Rn9sZpDbNvLRxGiwR9DDet7twaL54ud2801YeOfKoCcalXcHb1u8gV27ukvAX0o2
V5TgkyoOvPgS+4vqKOl5mtgtSibS1EB+tOPddPd27q8flfdQArfC5vx3K0otwjDfNEo4Ikap0IIH
kxND57Inecr/6B8rpnbjiBE+OZgSRWBeAFmUSSPvbseRR0VxfsVSgQHF1JeVm3wcOcM/5tH0eO+V
EFhi1n9vuMyqNICTyf7xnj8sSnzFiBoaFPxEZE5Rq81faV0leIbPYrt4KV2+PKLPIuzmThgcvbzO
Nr0O9mdi4Saha09Z5uAernGyd/SeyTkaEyX6MZFCHj5z1V1aKRjbp9eCcM25aGJL1k45FaaBcZev
cDGnIckUzKQKox691fMsx16EbQ1JP2xY6NmRA3cf2tnp+F7xchkUgacPEiTXjPAqv+MStBs/knU0
mc3Mp2RuJnNJIfTnjZlBd81xZOpCt/dMs5aGpfYr0fktUKBH/OyWgKYrleIHSNw1GETgT5k2dnNH
kn27NcxMJeu3cBuIxmOwjnzQGIoyg6I9Cdo68gs8yQLw8d0eIptDtvk4M9Jui9S5j0krkP0ddhZa
fEzUOoQa2nSgMUGKgnVife185/mmwrzYsJbR4/qDnWLCc9EQfIM8/D8rKthHK4F32QsN8ZfZ3OPM
3JpVSA7aLzzMqNVCGPnvh60BzKrtvnuZqG3KGJ+sUad9W/MVMg/R7s5eTQDquNS7oWLxg6U+/bbq
pTkw/WUrcoCvJKY7vGFj1QgR6aIhHv8Lt9FvYLzTjXw78l3pslYGQYyib7iy/7OfGfBUStOoeqMi
jyZ2UaGDQ9tjsGZipSv9k+d6iqNzHBPMRAWFBaeoml5Dg4URJzT7hhqEr/GagXNz8KXGCceEn0MM
3JIJd5bNsAL5K1G1p51fwtx9hrtVINNxIqRh8dQsrFgaTuUZFuDtQMaGWfW7SNiCyXWfTw6t+D/U
ifIPFGUVkGbort0QUvJdUevsEhWBwoi3C3JVnfy1LdFxfSrFCv0fDQKiqAEtJE506XcIeatro5uP
IqPgpKf49Effm8J3yTk7u9ekxPDUqUNbh2GvTBIFFXvsGs9X7TOJEmpTJCWIJyCEHo3QbdBOQMX1
IBvKviDdEGwYPffgfxg5m0d+axBoeWkhqGAjqRycegRgxFyBLG8wt6LgMciS2jDGAwLfKp+MK5EU
D8Js9wBJMEiZdZwn26+C5/jHW8Eq7mcDpveAjA6P3fz/mS5Z60CVlL58NRCschbgcE459ZvJx+NE
NFZDopg3bEKCtzZOx6vZb5S6vE39IoPjQh2aP2jIuvHyy3WojipzUJ4z4YBqMG1ZEeuSzzmxYMXD
Bf27NxycGByFpUk59QBU8geeX5vIXIgT0XUJIslXbY63HE3kG3ubltOD+1gJP4mwV0FZBmopJTZx
QUfJHvJeL9YJAxkCI/8dLx7TbSPp+JQAooCPdIbOFVA/Tr3cbVdbf5MygMiEuzgmx1mZCHaEoR34
+TC02v6vQUmLx6pi9ZatkWiL51rD2cuuKnsbQ6FsZrbhvYAtzVJMe4CBZ06Kp45/YF6BDG8/L/eF
TwFgarSUvDTuqc4siVBX6iveiWikjS8qmhjcYiUYFVrnnUHTGyEAPs2Mg+yYv7Xoq9GnRkdpFIrg
wq+OU+WhX2s2m3ncb4DyNFmyipqsSHanZg+Cb9RjUAP28daoDE4+wQGUSTAvD3cUSVpTU4yKJvEX
SNlNKcyPEQyjcH9u+/ywEylBEi50pCTGFzZ/LZF/4Q2YKIkt9E8djAPtnMKt9g04w1ZkUK9Q3M6i
5MAW0j09GNZWFharzmo2CVZ6S6/0a7qmgFp2/xOZi5XG/Y83+d/yt9kBkaV7cMr1zS3cUYxVM5kn
sHtahlDkV8y7e+3BweeMqfJAU3Y5KB9oaHCpvnSRfwGtf7vi7Y/tr6nlw9/Hlo1dQeryNAWc2xB+
NdqJJZGg79OuraQ7Tw2CVvaVCy2vbJXv3eKn0LFIuBAxCFN8D/44UwbYluIM8SGurEYLcnwDlQEg
0N/6oMaSReGyXlA26DrXJaaj2t0Gz5bLHIUh6hXH3ostChkb2eHZVjRPBJ4X1cbFjJOputB61EtY
9Rs+WWh6mspJSpjzSbhKdtSlwyD+SAIZj4f0KmfV7OaTASail6vnz8hG1HYds0YRfnR6MEdKiUo9
3s9symc4yeuuE+Vtpa6/2lzKDKNAxRFZdlNVQZxkwFlyU1vZiFOQDepibl5wjaoPOivHQz5NdYYY
gZbGp2niJBaSO7LuuZsRrMFOeqGVhrpB6PF00+9ZUBv8ayCHOAC9kHXwFS+P3urxYf3nyYM5kOnI
Nwh3cGE4/nSDkWWNX+nAyMf/tQacGcRlCJfq/GL2/6icWPIhwnBmobs/D5n8z5hAFl1sZgQedlXu
I7lBeVRX/5p+SdYVLpcNV6LWkVf13wtKLYETi7nrWZdDtNv6JFLG7qx1XL99RgepHMUePx11KGk0
kpRNnIL+1+mvT3hEPNvgxNLz0UyAmbmSDu2dAuK4QtfW0huYdEHH8efMWMi/atc5IMq1JCxyk8n8
y/G2c7gVYqECXiFkX0kPw7PBYRmeKQVuUEEVPltDrE9KNQm7peQ/mJlDn3kylhQymbtL8voEgvI3
w+E6kV5ElsAsXs8MEhEwENRMYguRhGu34tv0v42zMdF79dc5krW/k89igfXmsTHfZoqBksekBQvm
1gCcEB+S1LdQTZ9OaHKwPnW+6wS3bytXf+L1b96AbIs1aal32gUK7vyzcENaS8KbNOWq3AO4x4Ga
d9ETXw3mQVJXjs+v4R/dxWvVJUos7QBEGhhShIcFgJa0ZGrkCwGqM24tiNwU0gbAejJf25s+alT6
E3QO2Rq+wLJp0c6u5n80KRiOpDqKE5dcDMQbxmXqBrCOOshpWG8ZNZKZpT57Kro/X8C4d3kAkARX
azppiOdKFBf+7z/Q/MISQSYJW7HZsvvoFqQkT3Ec8hLvKUUee1Vpbl/Cwu3mL+3ihDl0LF0Y+P5w
dgo0s/I49d8ToHrEJKzfkrfOfziGUH7k8cPcxlxX1TlXT7CfEMwY9qNwcIGVDzekTPAse7/Mk1fu
U2yWa05ppS5qDYGN4Aie/j6ZO5fHD1hr14tX72gqmH1gUE1YfOu7xpp3O9fDvESOwsHtiqMlJZx9
zeZ+erK97b/qL+lPROQ7S0L4hEuoz7aQbpf92WeuXIX/Ddmnbc6KpmypI9j1w1U3FsTuT09h7Ml4
Qlu8oO0ueCekQlSpcIgmWY7kouIV0t6eX8wC7Zo4Efl8eZGsPiR1wCZJiWUcQ2R4HMDUWxBZL1QJ
W2Yf1RzDBgv4LntDKj5LCa/um+Y2nGEi0hz/u/5bbKuB5REEpmgX3hSUlhcCyrFS6WuwNsGrHKmA
jAF+MvycfDT7U55C1s0YkpP5G3m0Jwh/Ib1InlZKEy18ql1m6G507ALwYvgyG09iLvr/09/T2B8B
538s5IMgtby9mvfOPFquuafXOktSR9o6NZOicf+YEIYw5qF+aLvJ0s1kds7ipJkWLASfPr5qgYom
22LR8x/4itOaEt6d0MSS8X/sSnDiDKZLdeQ4/mF9mlvFKbuXABoWMJvJOwMjr+pkbO31ZsScXgsy
ZYV6g1HJXfksQUVV+YMIiUpwv1ztXN3LOb4lZ7V1ci0u+a4G2JvqT7QrxBMINxCZPdiuvQZthp3W
dRsKGCWrotnYFWotbLP100P9wCqoysDFrZ7nf3I6iRb10BAa5b5K24bdVMi0TMhFglsFAhuB7B5t
e2SmsiyfxrkQiGhgOUVIUBxsKHuNbY+/hRINlEKjmd5ozvGcUiLW9/58tXDTZ1yoSK/bRLBD/QjK
VyIZv7v54kvZtYVP3RDBkVk6rUxVn/tpPCrPd9FfUBMCXbbsGlJdKKlAdLGHJZ5gvHt07lyNqj8h
g0Ud3Li+CxXHlYM+95jdYtvZ+bFbQLGp6g5Dzf1L9EK9DP8+Tf5VGLW80w934fJXhJocqGkZ4Icu
BWaFisheXdKIUP8/lj9uhE4Ge2T51LMTL0Rm/PZ43UYl1gERbr9ZZwT0DaTSA5M1A9tC8Q500nFa
d9YoxNcHJqgDevzM4Xn5TN9vtyLyoiGS7MegPk/DE45XIl48vkRu6rGsuLHNZE3r5JoRcJ72+Zk6
0t42Tmd3MaUV17djYfHzX+TNmLNATgEjKzw7fy3oYbN1ZlrcHV04h288GQUxdUCJwqYhH9yw14Vj
ICY6WjCZ7XqSvvGvJq013QbQPr9EwSwneIGa8+yYN0O496MRqIkFTfZXfP/YprRPJaixceKmqAdO
Ru3u0rJVQSyVdq83c78KVfltc9oucju3pxVmCRLjShBzACNh/2TL0TELOHkcsKdyDKpvjrOKCp8c
tdMW+nShSSNBBv6XICZ6LDV8foDgaOHEQ0S2ef7k/BtlTIdhdYbQ8zJN5lBjFZ4MrEonTi4MxwPp
u3jp+xb4859hKpai6Ybegg1NTLtb1AY5cclDorww9liPwEDiaJ5okhOzEsXFsxZTBc+cyq3qRaXM
aLRpXB170d2+X2z5ActLD4/nJMepzpKlqGoIpF3dkBhNZr+tfc7xkNDsAXgA9dtCEFoRHmMI809z
9JVssN/ZWcsoe8sfdr2gHeYOkPTYxPQySwKkDmF4cAedWy91oLHxE7JYPQafrf7ngPx4VmWdbxcZ
fQyDsEcNwsr67z02kV1NYV8VrP5o5xmkxNV7xfL8Sq5prnrXw8Tw0lLRAwXgPdaFLgSUh3a1OK+p
Cxnsja/jMiG8D0F87dz2bA7f7GQubyvtf+zbxy8dh87CZEhnkjOdYNbwCDhc4jLUoUCNMYglKBml
YG++OHZ7xWvLy68dnEQSdGpojpihQMA8H/rpsbb/myJYcQzJ9vohgCn8PUuLKzmvvkXv8d6MCb0W
Ou8kFosS6t6Kz+3WBBilRlfeFWqNo4kYaCqsZG3UZs8bxpIwdkzPohmPcQPzyXmIH15M5ZU+HRjK
U4o3uPVpqQ45dknWSYMcJeC9JG9zIrFsPgu/kEuE6igFUYC0e0PV6A7NHzXEp1CoepkOMkgCKHCP
BdzydUzpmTxWvSI2ZuEA3Q+6iSwgvf1jCg28fnC1/fEziK58OkMxQPVT1MKsZi3O9yZbppbiH+Py
YOvBEOy3VYTLlDn5hEgSUavwoYzs3SSWpssPUe4ZjGIPkZdviaXr4XV+gDmNQoDlTZZSYkFoqB0C
/P9vFc3LkzUtfWd4VggTDlELsY42I55YfDAX2uS6WW2Pxrup3SbWymuNRynlvKxQZlZariumiZS0
Fj7//SBodFoFusU7c/3GfabC2tiwKhly+IVZ010Gl5xd/gzd0FlxZCct6jVzoa/7u1QLAGPo+jIK
hf/MtiQBAOQo+NUni/C4jLTBPAEtPq1r5XRVbIEnBaydifVOjcOhF1XTBuyeqx914ftOKGQ70UVA
UopqQ+FxT55ryMtIT8haEQcdKMLHI0NepJjOZMSre4Bh/jDpk1wBRWYiqb0IyzPtasvEWIfAmWmU
4IW53WWZytUFPmJuF9p2hFw23CosJVYljjRGh2v9EA77tPPVF1tpvvi+pnA0ZDj7a82D11REG2jt
8h92xmCdNqN5x59Pb8EzLweu+b7iqPunUGK20hp7EzTF+ucuG7zPVBIOItjXbVHS9xRH72WAXP0e
Gk5QDMKET8bXhc+Q9VShz02edbp++C7mX74i4pkGdvlBhVzLjRiMCz2nUHJ1+YemBGndBmBwawxn
9Aek08vEsUWfSynVoPGxt4mIXOdL27sf0jf7bO0RCAkFrVWFHciGWVWQNlsY8L7emLIfhYdwo6Gg
JRiKkGI0Vz5aNbMN9k7niknKtq952+DZ18z/0tQ0An8bN94Azn+r8JyGz2yPZBvYgLbY82OZLgAc
xenLxC3sXKrgyiMo0SSc/F+2webOWI4ygGAr4tuJCuC+yqmb9bvbH+bW8ak9PHOAOnorneD0kS+4
9J7/o7V22tp3G8dvPg9ZnR2Su06i0A+A+CoMWefe/oDSiPSiXhrn3Qjs4bDQdr6t+T5RJw5mBUd/
KxfVPBjOvjUv0EjbgNcOMz7xKw9qYfyWGsVIKamDL+3eS+0P1yoD7mkqyVc26IoUcmUWb3dJL+/V
u+RGYLPRq+GCx/s91Sg8jvrC90hgP22L1wf5I9JycP+9Ge/JNffD+FIq30aH4qR3ijlasICw+MVO
Qn3AZKC0yEVNdGZ4e2tLaPvm5HtP0csXsC2hgZ9EPKTwJpobjUvq2L74CsGVTyJLsOB1zoCkdqSn
EznWMo670AiV+3QbSR3pyUFhcFY8Dw==
`protect end_protected
