-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
LIuXXS7LxttXY2K2AMlXmtcSPg+2vOWreytwZKREYMgcT3cTpXzwezg04BEN09FHgx0UX0E4/IQU
5YFOV8uA1bpcuKecIFymZgN7kaXt6wbTGCNmbiAdGjIEWHJD0mE27P9uln+FGEA0kCEyuLcV2GZU
1I4VrRTDMR608IcFzfGBE2VZXHXcDJiSLHiOf4dFKMtFZTKnfhWqqxgKMp5CKZ9sBRZjHmgbxQJZ
irq8+nExOqPP59WuUw7CzamMdyptBcCMySDEDEjBc8i/KYwsOTMcJtiCDG2Tao1FxKXu8rEvbCpd
zki4HQnJpVW39dmUSi+/1lUzIDnvkjlUfMNzQA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 3040)
`protect data_block
gWyaFUydtQ/TWwOy1S4xsSE5EdpIYMDazfTs89/SJOZj71gVTbNumiXvANc7e+tm3L7ducniZj6O
BPJIh0WoJSk/tQPGD4EtHVRslnCkgW/8qL/HhAi/2VcJMFygPOXUvcx9QqgHJ8KkAJb+z6Y3vNBW
8MkTv380SKCAaU261882FQKarUnkBZEzPqu5nv31srvVDJLXQDFMQ7sDNQG85qOQhjCQAVxWDJPP
FL4ZhEGrgD51WdSMuIy7Vo66DZmgNJyRMOyiLhNm3tC6ZHxlb0khqS1kSom9Qz9y1qsEFd//6SVy
G2BU/nI4VvPFr7GmAytIi7HUwj3ykxdhYzLrUU4vzqUI2e3UIIMqdugck8kYPIOpxy3LMWDJ8BYD
coDAszHakqKnhGrvOd+zHFePTAmC1UzBh+cWduWYtkIZFsrc/4GbptiSl7tzBwWMQMJoua/HrvaH
X1ObF1uCFq/yw1pdwiBtsc/79McPeEdVSM0xyRstJI+t1qbXwkqkZ9ADKjManqr/L7Bh7B1F2TfY
l++hw1RuN/HmnKKzgYwyO4/2y3IXPDwIDBKdi8nS3SEOizjitlXyH6MBZ0+Dix8S00PrnBR40ZnL
/E7jh2zTTrj1ml+4nzECvN/dUjjNujXE7dLXg+U8CwlDrYC1jepaYQ+IaxmVOOfcISldeLh2pjqS
8qqVFmoPoyTA+K1Brbi8G07LAo66E699NSU7lqLCHUSMlbyxhqUGujOyRUpAgTlefj+Dsn/SpYir
5+MBJuwJhxxKsOjWBrRVDU10J8+tKX4bYIk+gKAuXk2u2+5Ls9yRiBj52WbBGrPzIJHOExXX8ZB9
iH0qzUfM74TmHhAjg4RJKb7G2PKsNQqKYfTAtZRa14XAy8X5q+GzDIifdR23ob+0t3LEcM3+FoLZ
nUQLJyiUU0JR3mGpldPpgAGSMunZqoadpzDqgamsUKK51KPkAFTkdUluRB7BGTsjmhUTqb8y/Si5
ng7hR8ESBczLU4ipnkIJl/FTcx2Z2NYOOR8TQIIAXL2XTO15FUmFTTQYcMgJTIIktXnTEmm3UsGB
otyzeOlBT5sWw4Nn7w9Zawm9Prrp1DFjKaT7PW3MOiGI+bC5s2iWwO27cHZL0RpvOp3gmxBcNHOf
m+Gvb+md5kgmFyPoZgzPFvs0ytVPSmAw6nL1wIkS2m3i7MKoqHcdM5CRwzdR53/c1J5tEAcl0PXO
5RdG10h9oYTFw9jC7rztch3d7XSPYX2EJpEdtZ58Ga3i3QNLS52gsZvsQjKW1T5wclXIrGgB/eIE
vmiYQxhZfZUBpf2IjW+tX/qr/JDrDkeexcHSSMu1bXR/Wse64fibqe8HZsOV4573xSC9Egx2Pp6G
3iPVgacWxFPHUIQZVuuGAnw8h0cJUyPWqcQmvmkurq9Yi+/kBjv/7Jq08hJaGkRHHbv2GTz7IZ8w
+dYFEXSw69cBqpkM/GycFZNET1+UkvBYx5XXx3kzrCX4eYJYhC5IOzRPoX8CVDCxh0Tu65WkKznK
ZAqDK4vASulzaU439T7wKMXZXpYMdWJ0+WlAQHMq9qVnMUFRK+VHq5y7rq5rCS2NWFAGjp5CmJ2x
1YKlvSMBvbm76k9dtGI6TCmOTwmWf1YSOTgW+N/X/imOCaIwvy8AvqpMzrmAcjP5RrsQKN9o4u8h
/WeRqMXRBbzUvCAmf+kh52510LZ8BJLoyjm1zUTN+wEPRPuN+2CFAokcgK92SghMnliEsNoCfXRT
lQy+cjdP1Uhjdjn6EKzUrPVDsu96dMHYZUfQ9Wyqlzb35S/zVb8zL1iRmo2EQyKc+Rt4tMZ/jCX9
/Vvrhy7ejMvMfmWGJPKRJ5MqvUQFtBXHlL/7+uUVJ/VLo8fxRAntZvHzn+kD/bNFFnnUoK9Ft5WP
wJEGglouvGiz9wKNYuihDPl996Yha/ODxnKqJxyP10Dc8F925CJMyqkC5IGxCGdntN+mp7acI9qM
KV6piVm4AFYN7v3fUuW6aSmjg79PpuDtg768ZuPmW4dRmCMDPtpSgJ9sMDhGCaLjX0MdjiukWJtF
m+A4ceAcFFw2BeB0D1x6G+/Fe5J+CYsGGO5avlx2xBeIkjaont+JShflu9+qTXXzsdGg2s5KljSG
xM/hrvwB5kl8ysu23c+XoIYYJufEiOlIWac+2wWxlOGfEqNIvPSE/m/5yFgSTzlsLaQ8d9mAUtGS
C3EDO+RVD0FNyVgsQIVpmyg5M2RoVIyPzWYXupqjj1nEVhl9+rX2O0IrwKv3Q9rnES2PPE5g3yyW
sEslpcTPhv5JznbVeKITXkf57JVHx95PACzJ9JYIN5lhXV7s4GW6HqRVeJtwDZXbXCKJWb7llIIJ
qoSc681HdyQNdxJVxukf05HQATevtw7b23FgmdzPtOITAomvKO0/ad5JpZMy3ZvFFFxfoh5YZ9Uq
Q5bFkw9vN7Trcpotf62IAzwE/IeZMe3ZoPb6G5mkd4SGgL9B1MeE+IgOwutptGz1exoumEmCESwh
JfDenx20Z4b6VhMCjspXN9mJup0O/5Vg4TTAkQEGmMU6NymuxA2jZRv4mYNaf8wIv0n57DLoqri3
OwpDiEoilsHLFxrZo9HrORp6GRg38e41WFLNZjisCCXeOMhGP3TmHXcP9oFON5gWI6An48IlX3RI
J8D3jZmRpoP8GxheSNScY5Vx6lvcAR0n5ZyRPnLjGlsSCvdxwuXnaSnrR+x6/vzFJ5yi1QP/QHll
QaDWiWwU/t+OyuxeRMHIPqJ7SUBtp6K2BkwuXB18ILBffDGXccyb1NrLgVHXctcK9bjYm+DuvdZy
eVruVqokTUFRywfCekGkS/s0TEaeFL4jpPnu0vw6DpAqnDWMPhJ3w7L0y3lP93AdPvtzdFXn/TAB
OQp5O5wduGQ5Ai8a7ELCKBLU5ejfiTW+56edKTxJLx9bm6VT4BTqQDTxenbSnO4cSgGVLlkiw/Io
2zXr/u1se2VSbWfxzi+m7YG34gHXHM77tgC/YCJ2GCDNlGOd1swgIuTvua1wqdCDji394qNp6kGb
muBWiSnKl6ajhs5QUpLPOkM/e9MR8qGAX2+Xg1Lv5xzAT0AZ8215IdvCLe4t8GoDWirogMpQzAL9
uVk/tSIBwIzohrVROS4KrRBlRC4enCCBi9xpWZ4UDnppuAHinXKowbHVRKT0TqaS5ewmcVr7t7Lt
5gWT23ol7R/PZYXmTOqUYCP+xoZmEa7CN/MSB5K35CHbqWka0Xi06WuPeFyG/FQd70s9hk+ceiyU
LFwR7Byr2sE9IA3auVon1D8geg2SZ9vRieBky90al+Xii5uxGCt5w56ZuRhlv3tWswJyJAK4loIs
QfoTPbRqdQCWVr+MtUTohrtPDLePliraY6HqZcum9liyf+e776lQqJYGq3vTjMhPkU9bCxlZ5wYw
FOT4Y5U4MN8GZz6J1TH34WNckZ4AlC33HcU0oL5E5s53GPaago3IA2R4do1hf2WvfkbewdIf4d7O
IAtEGbRlavHr0/Gzv+HKa7pkCIq0aWlbrqeHcy9WovzaEYIssKIFtBD7/NHE1dgYyKbJcQTukDQQ
opKn0t/wCS39q1y8RQ0i22onUsUBceE8mG3BIrBNyurpXedYcCJu04TxdYCRMRaWcse1MeD/3bxv
68Ecukzgw0hN4RCfsiCksSCbfIOClPJ2p+sLQ8kJjQfjh64xrgBejhMSZYYodzqwhmRhNdUBV6hI
TrfDyulK1jH1jz505RD88/9/4X9yFK5QZif6zDqbvGAVNLYbYov6rOTxW6ZdrKZMDZllocwIuA2V
Eukpv8jx5cpK4PvQKZoYN5ycRGBc1t7Bxve5+mNt8rUxA3Gu/I85O4Nrjva1f3UyOWZyx241uK4l
JFfKaSHi2QEmoUhlYQJK8KMBpjAEqK9LzsoihzfWFqKyMtnhAYvb6ZSbgL98SlbDMQnymHaknFft
IYw7HZ3O67AmRjJ9w/zvilk4eSLSM9Ajx2WsPDaGqHIeU6VT/9Estj9UCOtBmWICOdkmwQdC2WMD
jYiFGhOvNQAGbTdVv9nqXbi5OQ==
`protect end_protected
