��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o�(��	hM�j��o�6�'��RZ[c'�#�wZ�����Z?�3���E�H<�V1dݕ�N+=�c�
褬4�iE����_! ��M�9លie_S��J��`�I42%��d����XgV��;��v����.�Йt�M��D���
��OdW.����$���Ǵ
� 	J���z٠��&�f��$�MAmV�ԙe)���v�ead�=8��,�cRK+������s�v����,�I��-��}|.A��������b�ES���,�MYk"����t�)�i=�0�b����oB�|Va�Q=�oq�Ś����
z���ִ㓬��zL��2���=��bN��Z
�yE2i!��Ѻ}em/𔘉=4�ًn4��*t���j��Xd�5�$�}���&3M4�^�$����b�n�C����]�+�쑼�����
)�䏄f�r�/5��)�~���i��EQ�������X��@-����r�]�����`��v�!�z�X������Ipڶ��������d$���?~��_{3��iGf3WW�킺:�BE�=���v.R�;\�u~Ux��5���ae���-��LE"�q&-�m��F;�O�����7���)o�_ؖ�	U�����rT�FWeAR� Jz;���D.��A?VB�ߔ��R��ꆣ��ʘj�}�p���s�6-�sY-�$mN�l8*dg��D����W����Ξ��]�g��P�-�K�drQ�ȣ�͎M''���$�\��p!m4���s��KA�S[���H��,i��:;�V�6�\w�?���yY��UR��Gĉ/,=`╖O���^�/~�J)��{�����u�I7��4����:�#?)��롍m:�c#�F�^�0)�4H�?��S��1k��U6!̔FB)�6��߷�&��>�pn�Z���=Ξ�0� �D>�w���Ŋ_�	Ѹ=����a���7J���W]S�����!3��4���]� ��;;H�2�B�>�Ǥ�ʜ)�:�Ww��k�W7��=��zU(®-���b�q��f��F)L\�W{�C�p��z,�5���Gzd����X'"��D�<U\�5�+�횊&بZ��y^���v�@E	h����E8�N�P��G%й�^�L/��@B��9�>jK�lK���0�GTr�=Vܷ�k�Z�{�d֢�6(!�u�:nbt.3��	��^�4�Av�������>ҕD$�sj[��v��0�a!v�ȺP���7�O|�8�%�����b1E���6�1�2�:zG�AR��<< ���RU)��������]st��8U��PJ��W��*�3-�ɛ������~�p��v-����;��-̐��jʮ����{y.!�QtQ���VH��ů7	�5�zx�i*�"1H���$#�5_�?������;z����Z(��!ϩB��YSʃA�������i�Lt�yi��b�-���B����	,��v��5�M^��Q� �������s]1-�'���9�y)H�!�hF��"�BE���^��X@ �-�`�A^��?(����6&�.�m �C��n{�}����Ϳ�N'�5RK(�?先M���O\�d��o�ӭƧV�G""1�K��'��b"�\/�i��MoL(Ǖ�n	U�1��P]w�l�	'������w�XU�d�-<S4�k'�$���i���$��^p���e���T����ͧ�VeI'�ED+w]uV��b����y��f㨆�������d�4��!� `�4/�:B��X.¨��y�)�d=%���S�J,��f���C(�z? ���C1d�.�$��!�5�gI���Z6W�-8{�ԍC��})ȥ#$��\��l[|a���6�[����QTp]�oJ�9m�]��e54E`uD��*�`��k �c �:�7X� ����D�(�s83�
��Nnp�n�mÞea�	<�ذ�L�9�Y6��YC��A�q� i� k�aGb�hrc�x�B�W��0X'�	M⚶�M��I�44��$�@��ȥ��G��R�<d�ܡ�jh��U�~'L��2���4h _�Ka��"�G���v0��( ��g:���Fг��Z���\y�g����9*�e̊��J1#
� �hV���j#�Rjf�!MI�3�87���6�H�%���S6X6�@q�y��Hx�a��r���JH;�1�⅌s��#IH#�Y�T�YC��а�C<���.uN��Pw��#��C8f(��Nٕ�M�щ���- 6�1�o1���*���6�:L��:d �i
 h�QZa�f\��ꔝ�fd;:����o�xq�_g�Y���- �[��=�"���[�0]jH3u�ͦ'���)���/!Ab�rp�0��^AѤرi�o�*�r�sy�����8I�Λ����cNrؕs�X���c���dѻ��A���b�J���`z-`���h��-��>��Q��6��>����X��fa=jV���Q�E�%_�����]	5�t�	ȫ�;Z�1�ګ�|$۸@[O��S���}zvld�\Y�X�8�>�f-�j0^�H����5�RE=�����?��1D�yJX��%�G0I�  0E^f�D��'O��ypߚN���z��Ι��y����i㾖���uAk��Bƒ- 怋)H15�ӱYD䶶w0�ײRg&��D&�2�^S\;%����*��,��|I�ˢ�#���n78�+tĬ'A�%V^��|���2g@��Hr�7�Α�R�2�Pg�́�nn ����#�����KȈe=E>9�-a�n1���q@��|Zmn��������c����\u�Ԟ��m?�KD�������bb0�ү)�f�#�~MϜT�֛����Ӳ�'qV.ƚ5�6�|�`e��t�.���ἕ[�D��'��W?�� �ߧ��V`ޔ��L��
&���^����k���8�
/)�j[2���FW!��6کB�#�̮�r�F�60vtVR]���T��(��n�7[�0�+�X�Iy������cbѝ&��h\B&3$¨�w�]��~����V� ,�N���B\R�Yx���������h�e�l������mm���;B0���;��CY9�M_[�(7� E���u�j������Y؃�-�ւ5ʃ�����ʃ�{��d�7��Qx���֊dz����D���\��8x��a�e4��a ����!	�8x��s��9K���;]z���'�Q`.���<��?Gh�c�x�=C�vd�L6�E�:�D��~�C3�<m�ve�i8}��p�R���\n�o�
�9%������vz 9AW����5ƈ��6nwedY����� ���Ϻ�9��o�2���>m���z����E:�nE�Z-0�M��K�i����y���;�w�N���z��7ǟ�Kݿt�ւ�7˸u�����.�A�(M�o��R�k�quTK
����т��CZ_Wԝ�q�k�Ksu�9��KO�Ch-6*�N�H�jX���e��3�^�k`������e�gv:��:a�e~���7t�y�����6���ڛ�(:*��w<~�����*@i��8�K�8��qA��Hs��F����/����ae?��(�T�P�Of�٣��~�K���ϑ�E�ךj����;�Q�5�ڔf�����mY���>*}W���f�����[h"X?�/���`ΰ��W&-�C�@��~�-P�w���_�~�~��,���7t���@�eW���?���3�Ʌ�o�I����GE]��q$�4#?L$�l<N��/�X2�k�X8�!�6>M��X�k��o�m��:V�E�L�$��������y�c��}A����VS31��BSM���B��J����!�g+n��8�������	��+��0K�`]b ���v����_�q�� ��}�٭�~���Y�^M�~(BDKK�/�_�{q�b�$����@6���ϱ|��~��|.��5A�����3@>]�I7f�Bm��w*��*��)^�o��g��"�(: !�k���C[�d?�3+U$��!)sd�K��F��rBa���[x��܁g��k��/W��w`�Bm婘�J�	�Ή]�?)O�o��~Z�(O����˜�r]g��K����m}h;+�g�@��~�e�)�ـ!@8��̛P�Z'�v:�� ]�d������Z�2;W.Ё��Ғ���B���:n�;�(�d9���)��U���`�g�s��ܴc*tkDP�I:*6�}�W�D����\
�l��xd\�薎��V�P�(q��c))飻uT��o�Kh⢅7Z�2!!��%g�L�D��H��'ތ���0_���A��� =DSҩ�_y��R��T�p��ݙ�_�g��{�[T�w�G����y��r���V�0,��2:e�
ǁN&�qҵC��بjw~=�ܿяa�I��X̑+��qXo7���
��ΰc᳃6�uCHݸu+�s�XLrH�ѧ�G���p �zS�ɼ�4�/ 6���yf;N����d�V� �j}Ǽ鱺ME��2^��'��x�(,t��a���*/�F�����H���$������L�~�+�I[�é=���+A(��/�!�Z���W�^T�\�rN�����y'	U46�1���>v�X��g�1]��^wa��*��a����@/"!�T���8��c�����L`C{�t�:�l!������{0� -l�a����\��JD����B���;�=j��v�!��M"�@�?vAz����O�V�䷮H�y#��GM��_��#R:I�nTΜ}R!��6=Z]m4|�8ABC+� j�b؄�D)Y�3㰁)��|�y1�|��SZфD5����CD!���L�I���ԕ
��@�u�Aw�k��g:�U�3z��h�/���/Ɔ�<���r�!\�o��=�ᝁI�d�.�{h8�M>d��|v�K(6�8d�	�8�)w��%$xo��	�-4����}�{I
��h�����UM�k��T���v[b�gS�X@7��:x|�%�C��z �χ�ـ������ ��H����@�S����_��~s{����Q��8�t�1�ҖY��0�&��&�p���Kt��C�`�B�y�Z��+�S�(����=y�*/d�r�����6�u�sVJ�IY���C�2~�]L[�x���PR������g��}1��r�̊��=��J��.�� �R��"����N(e�"n�H$	Y�f��2��γ]��lU�:�_�Xv���Pm��A�zu�����v�4C���Y���,.[�d	�r�����mK�o���
y���R��$0�虋��t±༥�R爑.�l��2����4�7j>�<���9;՞���̳ʤ�.TN�Y�T%V����&N5��%���6����npq�0�61��Q �P5 'I7�*���g�g�2��A	6zyd=A�(L�D�w+Mf���Zފb��p-�OgZ.]��w�~	���R(�-�y��a��2��b��[5iO��f�l}�C��d�K��kC����ٸ� %6e�i�bFЫw��9���	��܇�@E���P���j��2�>~ӥ~�(9y���԰��� ��9�~k J���H�Ȥ \Q	&��K�V=���NiC��x
;yc����nE����6|���i�,H��x�r%F$��u|�v�ґ�lx�\!n�<Nim��BZfAh���#�9�J���\|;�d}H-V����Ism Q�����1��X�!���*atD���p��L��6���[�P�D�x����]B<_!��.�B:@�>Eۓs�����8�v��,{G�I���(���
�Y>"{�L�$��7�h���5���~�dul���2C�c��?��f�e�Iw��]�������6_���\�FB�đ��4�,�9JF���b�@���z�\}��=I�^�`dY2�x\ ��A� 3��kj:������U+qq��u0H��hA= ���+P��A��N�.j�r�t7?���dQ��[��'o��%�_"!���
�]��v���4�ٳ)'{��AM������m�AI�������֫ாv�{vw��9���ʼJ�GVU���T��F�0�{ͭ��2�y��a	���r���\٪Oί�: M�TN��{�����`��]��N/�&��� �u�5�D�<k�U�jҴ�1��{7G"}E�m�He��E����t=0�x��A3�%�����8r�Ν���U�}�hj�ax��ޑ�U�Z��gr'ܦx��$U���R��]�TGAu9��!����ZĬU���X�>[~!7M���k�(��ٛf��C�4}{�O��27?����C�#�����+b?U���ɪ���upb:�`t-������S�8��٘�֕����5���\�$q�h�n s#w�X~�������,����&
�a&�A��0�Vwnġ�p�B6����1K��l-�C���^����γ��4p��@��qz���ڒ�f���V󶨔��aI����۵���ކ)�!@�̀a�ӗ���tv.�Iv�T��*؍"�x�܊#$u5��K���%�]�7��+j;�G@���Oi�`���,/kw}eg�U-Q�hP X�v�L�3|,pH�ҬO�F1�s[�&	D+}��6|Iu�ţ�k�5��l�-�����+|ua��Ks��e!= �Dd��!�g$g��Ӻ;��7i*��~��0�rJ�N���A�?`��l�x�����	>�S�)��j�?��g������}ڑlz;�9�H�a��5$"�Y~9&(n�ȯ���΅�f�k�Uj���|�^��h.z�B���~e�X�>��ZJ�w�dtMk9_�;�{~�uՕ�{��d��^l'�:R'��,&+���(��S���t�A����½���+k��+i�g�:���~
[zPv�@�cp��t�@�9U*>�`,f��"%��I	�R��P�e���"F�K�]�ɇ�^����/.�\� z�dX�-x�8BP�-����n~� Nh��>\y5*\��Eݗ�ӡ�dJ N��[[��}l�lG�����tw�lmp
��8��*,-�d��<f���@P�����ܔ���cb�)���� 4�X~�L u��إc��i�X��w��_���Ŵ`��yDӇ� ��)�p��\ku��c�>f���ģ��j��ie���WU����(�Tܻ�}�0���<�}�^
�8��5"��u XP��(X�J�x2��]6}H2��-5!W�o�t���~���pI���xW�F�%ּ�>찀�;����ߎ�6��g`$�<kG�F�H>s�����Ԑ��\��w:_׬8-�]O�r��	��f%�w��y��"�1���R��(4���v�S�:N�^�C+�Oz��/Vs`��݅�W_?cVA]����Q�큍��b>��d�9�b���T���ZTL1J��Z�ZĴ$7�[PO�͑dC�CW�����j؋�!~-�h:�ح����nB�kF^(���`��UHT����x��]�a�
�ø�����(v���!����$=\��0�bM��[��ЛE�k��0��:��5<i7�o�c�m��!�Ҷ�~pȣ�^��㸩JDgL�{b�s�u��z� ��ר���zw\�7��8�� 6�[�x&t:�U �z��<���ѐ�`�B�z���^#��i-HcP�fNc1���xκ�W�wI�in�4��0�e�p� ��,n,�>��Ro]��G4����s���c�\���Qҁ.���ǝB>���9|�@�s����F��OT�/�%�9�N�V��	�R��}���@����ci@���D�GP�[�����O�T�XT.sP��-�)Z�8�������8u���-��<�����0c��c�v ����WO#�D��~jk}�g�X�l>L�IS�$�(Xqk�m�co�7�9.8L@�ݟ*���v?੾g��*��e5�˗����CEt�a�5�!=����ͳ��_]怷���.��V��n�Z���y�����q�p�\�ڧ��C���n�b+c�,9Ӣ�++KnuЛe�	�j(�p*���ੜ�͹૸��zP����nd�-�+�ܡ����2�#~�d:Jl��<,8��;ɹEǤ����k��c�K��Jð9g����Mild�|0��"G���I7���`����	a߱tQ�i?*�pMUi��s[ڽ�:Q�tj������5��1���=[_O!~�^�T�[	{��TLͷ�]��4�'ȑ���h	$����R�ybQ�h9z[e�y@�7Y�!@Q�c���y.}8�么�[T(G��%\g1�F]ڒ�q�/��MҲv4�U)_v��qr(�O�T�3_\X,]��.e��/�����|���2*�h ��X���3��q֬�oa��-�G:�%���9)DJ@I���8�B�>I7�5��>\+��Qb������#6_�C����ɽ�mQp�r
�ɥr^f�a�����7/�j�6$����Wփ��!�P�faw��1^J�=�h[0 _��!z�T��:=K��;�>�Z��u�!=��ע�G\BS!�	=���6O��mgedw�W��v������w��l��0�%��Y�e�%*}�
�ۺ'�|��]�B���U���'�{�������\7�qx֓��"��\G}�D�C�����b!���/��7a6p( �*��q����1��Y#�TO���Y9Qr‐�	�x�>�L�i����?pnW���%�p�����W{�[�޸��R��ЁRA��u�"��jI�֪�>�EV���D	)��8�1Zc���XT���ʹׯ�=���В����z�Nv�Pay�)(�P\��������;&3�={$���X-���!�L>�

�+�iVr�"���{'�\���@�D�HJ�,�����6���zP	A�����m>�G�=�"P?����As��!U�O �*��q;~���\6[��g%����]3!\�nٓ�������z	.ZM}Ş:l��8'�����6�ET�2�U@ՓޫJ�"r�XB~�y�>��U��g</�a�4	/+�1ЄU87����/CR����@r97�����.���y'`�eW�x��W����!O��_���P�͞�5�T�ʠ� ��q��='�W�����h��s��(�0Tua5�~+�����лT���<f��ⶌ��&�Q��K�� $�Z�S���Aq4��?����Ңiߌ��8��:O�i��N`���H���4�[��ojá��;/�:��������gk�x���e���=T�CQp���� �}G�2&#��q���z��bv�t�����1���,�`}�f�j���S�;֘� ��n M�����7�}<k�DH���3�I���R�*ϗ�
�o���k�O�0�	�7�Z�mU�&_��&��y����G���.���6k�M�5��Ar�Dڊ[��U�"xlc��;���>m��˚[Yr`U�)�� ��;=$r<�L����V��D�2�}�zN��3���x$~ޝP<Z�i�o��}��d5���6�)�`�'�4<�`vB;����k�h�+Ӑ!�*����ekg^��=F��X�71���}q$��< �`�ؠ����l)֚$G>7@��	����n��5����2������O5�n0"Q'��)��R`���;�0�u�Z��*S[OC=/\?]����{r�>�g,Vo�W���.+XC��5�<o"�:��F?�8�A�ݡ�߶7�Lok|y�3%e�oɕ~kX]m�6i8��~8"t��O�r{ ��I���AZD�j*����Z[ۖ��=�̰^(͐@k0!�o����	�~~,ToJ�>ėz��ͬ8r��8C�@gǊ�M ���}��8��n��w$��+��8P����?vU������e�ň��8ߚ����wn��)�"D14�H9��W3��DV"]s��7{�ªv�a5������*���G��M��8
G"M6�N�xx:�^+>�^��>��p�Td���[4�S�&ԶsNk�W�[�3��Q�rg�8*H"K���������5�z� �.��.DS�1g��ß-;1����t�TP���eQ���J�W��M�`��[Yre������R֗����Tۂ�Ҫ�����zT��U���5T���t�H;�F�"��/r�=v�Y�{'!X,{mD2'�b�����b9
-Hoӧ���l6��� .��W,���i*2��ng=R1� &��<�[}�{GR�����q��ナo�����A�"�/ރ����8���f��QO�@/4��_ǋ�Gs�䂁�	��6yC��>�����n@����YA!��,���#GL�A2��'���B����®V�ݣfƌ�m_k�zD�tچeX�$�7�:Utf��1���͑��.Q����ѣI�CH/+L��X���O�/�K����cT��r,R�8Z�Q�J��{z�RB�G��//�΄/\?
��N���`���V!��
DQ�j�;�+n<�kSȝ-Φ�WS��_���|wb�W|b�ר| v��(��Ԡ�?��◸e��55w�V�f\�#�5S�Ũ�S��k��G=�_�?�������a�� Q%�y!���FZx3�Ӻ� `9�A�'��Q���mkVZ��w�W5xj�n�l��9��0���抒�=���8��3"f�g�U���2��(
��͸��PUb�m\j�4çH)��
M=2�N:b��i�AR�`A2��l�� j$�'�P��m�^��U5��lM4�e� X_��o=7��-�1������O]ڔSC�f��a%��ʐ�����n�|?O���B����i-�W�q�O��DtwoSw��xl=�2q#,KGf9CkϢ��|߁����QB��oK( 	����en���d�n.�%&��-�P�rJ��*���j#���zTz�B
y(�XS�F\/J	�E<ѓr}1�k�T⟷�mM� Y�K��O,�Z���P����-�wŵ+*�)���̖Y_T8��C�Q�8��Oj�̖��;�|\�+��\�N�W>m�#K�v�S�n�+�(9W��V���,�>T��G���* ��F4�ޕL��#�Ӊ%Ĵ=�R�3���v2��ι
~3~M��Uq���!Z�@������ͱ
U�,�X\������Bc/�+��JMHxkNigq*���n��P[V��q�y�=g�a��l1����� ��G�o�D�猁j׋S�
/�i��,c�p�i�;��)-(%���A1����}��1u[��uS��wy�:%���C&��x�1��Y�x<e-�XW�S�->K��C�r�Q5�A���2-,����s�w,�$~���_b:�'�h�2h� ~hJk�(|�J��[�ƾB��l�Q���AՐ.Q����~��@�b�>��L��Y�DFVb����r0$�������=�yX�Ӽ>p2O�ᴀ�߬Z���6���%QzW��/��=�ek����%��,��_uL8��%$p��tP
]���[U`�Ґ{�υX(��Vƾ�!T�!Rb 4�Z�Pdдj�x1�A�9���40ɍ���?���*����D�(�Ry@�m���]�i}uݤ�iY�'ys���GP0�Դ5� ����ŗ��p'��dt�^�a��Z��A��$�zL9`9��}༥�fP�D4P�w	�k��xz/��5\B��l�2X /�4�����b˖ H�ڂu��M��_�~[b�Ɋ��o�a��TF���xG�}�,\1z�:U��;.]7�;Dۀ&��c�a�N
�^e�s	~;An��V�pR!�`����fZ��557pvA��D�85��p&z�.��-U|{n�xp[�f�Cڑ�K,���mFe������QCҨ߿
���
p|�pB�p��6�L����`�C#]���0ѕ�Lrό�����kQŞA7O1�J�܍�Z{aGCh�.f����J������)����6
�,D��I��%l(��P���(x�O����x���Ǣ�*S"z?��z���R[79�☛��P"�?<\ܫ�B�xL�
�F�XB�B+p�M��̻Ꙕf�C�s,^�5b�>��vῴ���.U;���J�}`:'�z��e���P�Y�땼�X�2��������N�I[��!C�	]H�a�ɇ �bX�'���*�iԎl�b=�{��Y��:5����o@�����Q|�ͤ���m�Pkt��*4�2�b�i�6��������s���ϾLD�j��_|/^f,�[f����z��0���ǅ�uS���q�'V�N�
0�l�=AuB|���Լ*�,k�r�`�{8	{w�C����6��"=@uŦ	��=Z��B�w�Tʂ��+U}LJ���h:Tj<��C��k���nydv�q�ڙ����5H�x�)��?�1�;�R�ux�"'�Jt��_�d��Z�2�h�U�e�V�{��8梴�Q4���
�S-�ųG�5!Fj��	�j��g:3���t@�[�
���cM"���#%��	�i�Xb@?�h0�=hwn��¹�_O[w��u믾_>��C�M�7��f`���&��b��|���z0hk�)��[�<�m������>���ltڊv��dH"!J%���._0Jxq��,ө�B���5��Q�O�A&�]Ǯ�?l�� i�\l�ozUX���֮yJ��A�ޓE��|E8\V�:��KM!EO>�iJ[���r��p�#��4
��G���QS���[��`cnÞ$�����O�1�5���ݶqk��z(>�ҧ�2��N�<C���3H����'����O�>z�i{G�E@%$�, ~�=[<9:y7���,NI�A��m��\&w8�iAFD��׍��������~���T���[��n1k�4�V}��b��2����֘�ݍ̪���;�d:��<cnW���k��cZ��ڋC�ۄ���C0�'��V���؄9B��l��wIc��RI��L���[4�����4� F�H�F���
=��_݅��d��Ϟ�"T�b_�U�t)�P�b2����cI�UFo�/�p�w��G���v�,B�H[`A�gs��+�ɛ��9�U��3W��e��BC�����R��U��(c�/I� ��a�dY�MAfU�T�6|��@܍<"9���u#	!����θ���ge�H�d#���~�]�-��S��sS#Ў\���C[�i�#პ��z�=��]n�bR�f�+2r��;�G$3`<ޗ���R�J�ͱ�oWt }����߭K�*��sA���q��&�11D-~�HK9�k!�\@.����Pg����q�+	�E�.�L��ަ��5�c&�3���A@sS�<&�xag�;�Ov3̅��-5�$&[|���h������>C���@�0���b,�C����/(H���C*R�f�Xh�=|�t��Y��X��mL�3�	��"�wF9��&x��R�ƅk��H �y}m^@hN~?�M㎈���4��B���x��c��eٲ�[m=
������ͪITHk}�MMZ���z޽�P�9�g}g[��=�n�%1���D��S�=�q�U\��AOC^K�*R���+U g63���*�+��O��=6.S[#`�'�_iE9�J��c��%C,G�Jr��z��:�L�-Q�FH�V,>�޶y�e�! ���R�}xF�Q�舃f��e �Ϧ��祢O�6h�b��tꂘ���U�M�b����8�Ӳ^��}�B@,7�2���m�]!�A��Ik\�^f8�\��'G:vXG��I�4j��� U m�ѣg�%6|��zz�k�G;�	C	�W�L_ew\Q�\���(��"pB�6B�v�z�KZB��p�ï"%���%��)�|xħ�?^b	���T���J�+���H	%�YC���q�S7��VD��^X��Lů-vaQ�uv�ZlG�'3�'�7��)C*��R�)���;p�"w�})���/��E�i��h(��
�P-q�aam�]�e?}k���(׫�{%������v;E��W���-7���J2��eЇCԵ)!���?Y��Q�,��Q�z	A�pHڊهB.��uXC�f҂�z����8�i'�m(��'�8=6Jb8��	�wb2>.�X%�9����lb�DA�{� y�V<�*X*�*�e�n�a,I�5�@��4�:�.-���f�V��c6�0�V�,���\�1�W3Q[���ً3W_�w��5h#;���?�_o�,$���3 *Ƅ�nc��nUTh ��w9�J�۱3,,x�=U������J��Eq�%���#q��m�ҾP�@/�
LB�Z�;���֕���ϵ�ڛ�v�	\jųKz��|���J;�Ʀ�[c��N�9�6���QJ����-}����i2��O\�v٫���-ǟ�%�=��!G#G3G�-OČ��߁��9��׃�?M ��X��@��D������;+ؤԦ�<1���՛+����~�3��aq���qDY�gO8Ԥm/�+���@7οX8#�Υ�`��N6��f��xE""��.P�z.t��<�r2�Ğ�S�X,V�,ЕzÞYZ �bc�
n��C*)� �� ��U�����h;���z�A0/�k���F�!���ˋe$2�MxC�d^8�!�[4�Z��Y>A���)�<� ��4�	�9��-"�U� Yq��\���;<�A[��E�>W\�S����R�/��M��ފe��K�V���@ ��eץ��LcX�L���q�Z��4ؚ�1�ʓ�(檫�C7FM}s���g�'��w&��h��x>�EGs< ;?��z9e�Ձl[�!�Q�W�5f��P{Μ����l~ݷe�H�jき7�YFc��w~{���x�ڱ(ޭRQ�� �6�q�A/C�Z��J��29T�t�y�}������n@�B��ׅ�+��M�gݷ�D��c����\@"���ʀQ<�� �͜$>�Iyv{��DY�ΉQ���s�n�Hn2B��ߑ���p��M�;�%qlj�M�ήo������}�vO�Y28��8_��@]��3����1�s�2G��(��u}
��b=���{�q�yq����d̙*M,�1���V�v��Q�3�z���|f&�E�)��@���{)�jJ~O�0oH?W�'Vi֌��+��3�{�tP���0�Rhɠ!�c*�B=��̠�7��ڋ1G��\}ȄvjQh�X�uT�(B���l���"��A�^4�ЍR;�bQ���C�Q�y���[�wo�`�k87g��~_i���Lz��Y�w��m~NOP�\xm��1��<��N�/��f8f�/�)CU�6��g��LO�a2��=����*�r�%+�-�%���)H����Ӻ�����Ŷo$�ij�`R<��B�?0������28��B�9|��Ǆ��G����!=��+ຕ	�D勊��]��z3������{����(k�F����o#	�l.B%�E���l�L��y�A?|\�"���
Z~��M���̻.����AC�\�e1��8�߿Z݀���^�!aݫ�.u�f�o:�Z��(;���mR��3��n���ya������a#��l�J�DU�3/�z!N���)#h�ӣb�UᓇR3}���U�������!��$�ג��Mw{ݑ��s,��j-W�;z �1��3�l��$�,���L5*o�G
�v;���i�.c��v�;��$P/�� Ŷ-(m`���\o�&�۳Fi���@��['0��!�y��5���FV�����
w$�Y�'�C���3K������w�J�R�bFt{15	q��r*��z-���⃤��Lh�����Bv�gt���!�*�O��7�aW7�'"^N���n�.�O����Q<�Jv�� ���+��N��CH�Pp[O��k.�H�{��"������\-|�;�w�"��w��iS�n�ѩ
�&�������s�1�)�H�uR�xL���d�\Ix[�(�`�:�b������v�~B����8	�:��b'��q V��+�C��t?d!&hs�Nޑ� {�����m��r��t�����b��
o�)s�[��g�D�Ŷ'�%O��r[�l��DL�E���60k+�m�hS�������|S��t����"N�����1(�fcJ�-�ɺ<�GQ��;o3��������Pyt�N��'�	=v���(���BnE,I�1�P=���-�h[�� ��� ��]�u��o�I�\܅�~��
��,��ҟ���wB���vVA�='���!#�1��/�a֢+���,�~�K�"���y�manE�ް��?�˘3vFa��ŷ�<���|���:�S�*�)�&uhAx��q��|ÈB���O�{�wgm�\Ǻ �� =����xJ�V��Ԡ#�
�?�����`bLr�k�;��귥�h�Hx=�_Fɀ �9t�-�2u�c*N�L�ML< ���\�+��4�P�,zi� {N�{r4���7��^�����p��O�jG���iO{Y�0��=�Ybb`l���6�%_�ߤ��8!������w��L�Z��@L/�g)�y���Ʃ�wmX��A^*�>f	��.�-�H\�1Ů���.�W��,�1x�i��n�o�"kWW[��g��L�(�Xr��b�	�4+�y����N�#(Ty�<��#��l�"@�?�`L��P�1Z�!�+��帉�
�Y��(g��o��h��[����s��i��ƣ����R&+N���t!�	���� ��w�](����w�3�>E�+|D��I�B�׽9|���o�P��ߧ&������j�?��D����b��i�	Q�%��b���L)S~�����BfKB������p�ųZ�#Qe���4D�{��=��@볕�]H�.�ERf��썕�V�Zv�����k��y��e�5��u9=��+k,����b�h�)"��3����n�[l�;�_����uh�Ӯg7D%��W� �t0j����X��M�*>_�W�Y��o,/J�}ߚ�<�R f�&�M;�	ş)>]����45�L�[��?,?�q�U��Ώ�Þ�(�@Ø���vA��52E�S�f:��O0ϲ54� _�1o�H+F���o�͹�yC
��-��+v�d��9����^���xᙷ�G���%�m!*W;�]���%��3��~���^G"��՚���]&�$��:�K_���H^�X��aPT��F-�y�a|��ӷ^���WW��g-<������p�~R M�=��	�6c6�y��c:�~*��M"D�[ ��mm���0U�$XU5��z�3��7�hxH�U��[)���o_��3���e3B��R�MoX6��6"D����N���Z��%�X��r�"�"����UTS"���-\�7��/K����
�A�X�����ހ�8Z�
�ٙW����� o;�-c�ut�����c����q(���n��K��T�U�
�~�u�3��@�?fMqW�������^��=t΍�h ]𾏍�Gg���Ò"��\���չc�罗G��}PZCJmh`��X�Ea�h�!�Rn�]���V�5�ɤ��f�V�ʫ�5
��W��"�V��}4	,'%��wO��_%��1��O ��Z$)�NԷfޞ	mE�0'��$�K3�ͥ��a�z"�:
�3��~s������y�!����T@�uQ'�O����֛��F=�3�gaY�s�f<�� _�-z`B~E`��Cɿ��1�J�Dd�a Vb7�V�Ww��x�Y�~ǯ�����@����?�<�f�Lb�)C�7���~��/���kN[&�+��`o��q%L��3#��p�	OЬ������;
'�n��f�-��j�k%����B?����\L��U&pe�ә�� �����37z���6U����׀�Э�ۍN�R*��i����){;�5�BA����#�_b{�ӭU�!~od��=X����g.��m#B��O{�����S��:���
���� �Bd�g��D�X������Mw#��(Bo};5���p!�'1{n�q��!���OHb�[o.x+�Fqm'�xI|e����~k��n��Ά{��E��w�)"EAѯ���\e�PS2뙤R�WkoJX�Y�
�0J�M#��/6��$9g��x��?����ͩ{�PE�x�p�p�)��eL�N�H͟��ĿaEr�Ú������QweZl�RQiBz���(R��s��S'�y�����R�F�~YO�ϽED=wt�4��k
��A�ௌ�%Zt�wW�rn�5D��n�Q#�Լގ���]:H+0�����P�s8�+k���ؼx�ʪ�'G3�����sK�7,���c���ˍ�K�o��:�F6Ί���}{��:�g7e�:����e����ݘ��'�[�sq�]�$4S\�ک�����}]LH먯��{�E�����EX���l�C��~����MP�S�1�zOo���� 5YL��N ?�nj��K��/�t õ�d(W�"T������۫�l/Ƴ��v������[�-.��3d�Ԗ���W3$���臬i8F��x����_��R�{Ƭ�_��n�tŁ~���WV��6S�Y'E����@dHȬ����G�Y�.S%������G����MhR��`e��A躦��LR���$�5*:rH�(�.�o'a%���䩨�L�W�]�B<ښ>�����V�����L#^�c��H��ܓ޷oj���h�.��kDx�߫�F��~��.�b�hRj�䥺�Aps�+;aN�f�.�*������vx�T(�M����]�j�
u�+�c\#2�}�(
��7:}&�ծP��`�3�����>*�g���P��?�* �h>OE��~LͭU@�9`c�VU���{k�F�b��e�+�ķGo��w��?�^.��*���Z��L�~����T��?���̖�}tnI�)�C��4��!b~�D��B��
ʊ��ض��ϡ��qB#>b*��$M�7�#e���.-s��lփ�Z,�ݏcÀr�E֢Б( ˌ����\�~[�@3@1Į�|qn���^���3#�Iu��WG�t�f{hv�nK`�9&���S�sO��!��G��:w��n�^�9lhtٸ��^qjk�,�4(q6tI����Ts�|O6��ɢ�ɩ���|[�_di�s����8`�4t^_#�:!=�E\����=�Yb*n�.O�~�(Y�&�����-ϗ��[t�b�ڙG�BT� !bY|"}� ��V��]f��v;{����h���ܻ���P�p�e�w32B�x�uU ��akO��#P��'�a��6-GS)����t��M 9"'����t�Y~jgq� 2�����ۈӳ�	o���WJ[�ߠ�EV�]\c,�c�񊮇�u	1��M6 ϋ�0�b��0,������
�҃�
D"n�m|�7wH*�B����4�	�N,�����m� �\��ʜ���!��'��F<�d"����o�%ņ��!�j���B��i�^�L�%��r��܆Q�ӭ@�:���+A`p\���C�X�@4mqJ���l��w�_��Jb��*�'����4��c��$ť�Z�t�!���0}Ņ��21�H��C<��U�������ש�7�|�~q��P�6�Ϗ�S$�l#<�}����`�\�\H��ݰ��˸���0u-����B��K�֐w�A�T��ٱrs��c�8;��eS�� U��G��n���Ĉq4����ʑ����n%����K+:��h��[���S��k��c�Vk����q�J�M�S]��c쥬��0�����D�� �=Q���!�v��%�4V剖TJ՗-b���ǙbQ���7{K�Fީ�,#�@j�������{*�۷��Ÿ���n�����Γ�P���(�P�.q�%Y�jX�u�CV�,o�ZG)-ڔ��|CJj��Lb�<x�|������P�L���`�TQ��W�����ƪ��`�:�n;�Ɲ�^��W�3��Qp���A������]�����B���d]�dcq3~�`v��6�·��Mf�w�z����p]I��	fԩ-d��#�T�h
���ف�����kl�g���rCO�4bq��LR>RX�Vk.̠��l�����V�J���y�pM��Z��^�D����V�wӓ%�ܳ]��b#��Bs����T@�?ig_���ɖ��&���{��S�'�+�J��y�$4�� r$�����P*|{�53��7�7��W���9��F kS�:�H�M�I����ݹ!�L�6z����Ad�z7�%�z  =׀�D��}���)�0OP�I�&њ��?sE���-�> �-8��[:����l�Ǽ�6K�MԺK�<�&OUr:~G�vME%ѱ`@��� �)GV�A��\��f��ER��fc�u�k���l���ΓX*��B]�@a��X]�X�9�]��#[�߇�i�/����3�*zN�� �Y�뻪8���V��y�g��Z^\P/��E\�0	B�:*OcKU_-Ԃ��(\��6��Q�TH\���L?�uGEҔq�{��!���+П�/M7��g*&�ú!��f"�np�o'�"5���\��E�͊�ɽ��6�ˍ=���4��W�u%'j[J��hb��,��+nV����l�N@�o�Z����/���~ �!�}Sk����?gf�`zC�:b�G�W}�w��;<m\�sÓ`K�~���.���F�����������o���w�������+�Y!�:��M���M#L��}�����v;hMl��{���I�B�2���NX��*�X"����d�k��V�c���x���W������L\��=R�FB�����a>�j�n�ؽzW
���~-���j+ݰ�R�D����U+��k^�����M!�}w)"q�G�i/5�Q�E��_�V?��y�i��\6����4B����uY��W�,���ꠎ����P&���
SIR�"���޷�S�%�!�M��Jz0�k�
��&��+�ϣ
�˗�0(j���T�4�}�I�!�_1�,�`c@�]�&�J�ڟ�5�u�,��"��ߊ� �����ܢ��E�&�.�DP��f�m�Ϡ&)��(D��Ytq#Z�,����ٜ��n�5B�WgV�ȫ�;�0@Jd) �e��E���E�$�ő���I���c��c>���ŷ�m(qR�7��ZLC�Wet�.o;&7yO�vU�c�笆A���yl�}<!t;��4c�����������Z������0> =DP�$�f׬�z�����Ȋ���y;.s����C��\��j�:&ke_Ɯ�F��jU�{F��^�A+N@��oٙc����������qѕ�[�5}y>�(H5�d��3q�"�ۓ��J|c�ID�r���#G�G㽤w�� �>�s��!�y�u��[����l�[�c�;������*��)l��G��7�#��6�q|�@�<�[���r653*�K�3���@�3y�zr�)�u��+r��ƿ贇�
��T
�l*�㽼����B�T���Z�]�9q;�6����� ��G{J�LҲ����w��C]_�ǱlLf�"�g���H�`��{�۪$�+ϒvHBHA�6~�!�yf��������� ����WQ��aC7�EgT���~[L�P9̠u4AS�H9I(K0���A��8-}F�A	�f��K@E�ɐ�)�Mt�/AN���6s�sm��V=	Ư����X�0X�y�Eh��L*{fqAe�sl��Μ��y4�hf)N>F���?�Yv�j^[[K�=��~��$��������Qf0Sކ��L������-k���'O�f��{@�^B��]0P^&���ds>������~54�� ���T����͏sR-4yp�fqXz'uC$��b[�)�>�V3q=9磧�A� n���.�A��C���1�6�8�ö=@� 1�l/~�^6�)��5��?E���U��N�'�x�\Cx�<m�Õ��m�,a�^^Ƅq��*3+���F�&{�|��u�� W���s�_~������/Y�p"f���N��?� &����
5�K�K�$x[�f��w���
�����J?^�[�����"E�E��{ǃT�@�����&��"b���T�Zӻ�4�e���Ph M�"�M��E@�.:;�`%b�=�x�P�iί�3	�'97�k�4x�n���c��ꌐ���2Wd�Z��Ě��}��P5����:�l�*�)��Ħ@}������hsw~=�}uu�߂	<�$���h����#��FMVy�y`���ܹJB�-���q%�e֩�����`�ċs����@�G�{�]YS?�c�̐��f�
��=�5��c��,�/3s��c���Ӊ{��Me֊�Y�7*�MI{SoGx�XJ��}#fq{�����V��H�5_rL�>� ���_ɇ寐���#��۹���G�O�F�|���J���5'�����/O���	z��]e{k�QdS�ߔOw�
���G�:��@s횧����"�����*@���(y�8V��Tě3��xx���K)�$�s�W<�&�#��m&SĘ�0�����f�/��ӏ��'����
�k�g-���9��(I�V-�Vp>iF��kf��&�lK� ��4���e41�6�r?�Ex�����c����}�H�1$�@2Ù�(�� ����w��CXX����B�C��g{�-e���r�fJ��>�00hN��]��_���ʔ��L�����	\�x6�㒟|.���`Iv�H�g�Bx�B<++�Քg8��I�Ro����-����U)�|�3����t�����|��ǀ�{U������7�xȚ�9w$��W4褁�x��
�b��t�����z��ǁ�����	�<:�|������$0'	���o�߅�ĺ���w�g�T�����ۡ��L�I%����hm�m�mC�a;m�?�eɯF7����~����c�#���������g���`'�1�tH�JUR�XKjw�Gr#Ó�l��<��N��,Ӈ�О�B��sɮ��Y ��I��q��h�U��B������Z����j�,�<G,)�Z�걇�6?�_�w ��~�q�z���,��M7�A�l�Dn�yNd��;w
������>��h��4��(Y�������*����f1�ˋHZ۫�&N�J�z2�YW�k��<WhoB|̫�$2@ l���	.h��q,���"�Q�x�M�7eL�A*��7N+�
��`;<"L�JЩ�Zɕ[�78�`]��Y�� 7\O=*���N�6�#(q�n�]ފ�1`���HC��� �Ar�CTh&`�m�a!��J��fя�r&��ę�P ��4V�ߚމ���%On$���>��đpRT@S�B#�.oW3��v�4�dq�xE�8���&����P���²y�I@�ϗ5�E�|��f�/<.qA̘UT@>�C^�UN�抈��0�}~N�������0���En��%��Uk\a�hͲi��c����^��d8�R�Ӑ��_��ľ��u��\�4��lt���gr���F��%Ҥ,�ߪL�[����1�Ju>.�:糧�06�R#A}%����;s��L����H{�0����Qi=T�f�a O�����謸��٠��=���<|t��:ZۮP#�G�O��W�a��0Z�P��`�G9�KR�-�_�n�6��0�#Ls�ip�f������|ڋ�R�oW2e�� ����쾉	���#�偀�������K�7{�5>*�Tb�f7�g?) /��o4�=Z�˨����:U|��ۈ%w]=K'�
j��|��a�=��q켺y@|���>s�Vc6��"J���x{pO�U�:����[^ʯS�BY!����w�P"/���:�n�l�������?�S��G�����a�6�*������b�0iʈ��QEŷ��N�\�A?�N�X��� I2j*S���oE������pP�:KI�15dy9�^��[�ć�.-��;'�Q�_�6ל1����ҝ�pX�z��ϳ.�ۣ�Ë{�rB�Q��vj>d@f�=�Sv��c=Ļ�pjk�1	�d�ӽ#��c?Җ[ݲkȻ���a+�y˦��g�97?t/X�$Q���&��J��!�ޭ\�������w�
��S9�V	/atD�l�K�eȩ�`iĳQVVE��x�|���v�}s
�Ed��nñ����~������rO�Ys�G{��(�+�����V�Y�z0��2H��8f���4�Z��[>�I��$��XS���9�qY����ۡ�{�aoJ8:[u��~p�L����[�s�.u.�:�T�نP�4���t�|�Ϝn"[i��$�+����GO�Hc$���C�&V�:�X�i�I��Tes�f���D��H�T�����=\s��BTߝ=�;���`M�8����I��zߠ�\¬��H������]�G _�ۛ�u��׊䳓yG���ur� V���k�7;���4��Źr�Ry8w�\ES��%����/D����?�C1��U�z �\kBȝ�;]f�g�PȠ��v��!V�v���%3���]m�"�EI�"�t͕�)-��M�8o ��
t������n^�f��� }�JB���|�GѹK7�"��"���s�a�>�^��i�����|`���#�|~G,G�]��A�L��&�+��ͨF�+f�ٻ�9qڇ5��|JnL ��m%�9I��|��[�{^)�OV�3�~�gב�n%���u8��Dk����uҌ5W9p�+W�m��z��( ��Z�κ9E�9V4-�_���[
ٔ3p�w��-��W��X�)���|+�!<��<a��B��-Q��t	{�F�&1����I�=�[=�Q�A�$�8�h�G:9�(_E��{ĺ�L�l���t�t�[7��H=ɶ�y���5�߸ d�$�%yM'^���r U�A�O�Vp�szQ�~�[�3��Xk����>;�-j:s0�Q� ��6�ԓ�аm��)g����ѯP��|�Q&�	�%�L��%�D��\�k��2��_��M��A���fh,��}F�a�'&���&o�;G�k5ݠ�U��ꪰ���^(��,~�~���ěN�i�e�p����/U%���t;���T0�L��k�Obn%��<�p�pw�6ܷe��=�bz_�]=h負^�>�W���)᭓B�h�S�!��c��<1�Og�N	�hpF�DvYڱĕH�	=����y���zV�2Z���GI���w�R�ɢn��׾��Q���]��ַT�&D޽ɚ:�a%Ӷ�� �e~c��R�����(- ?�~�B�^Z�@ρ5#0���#a|M�2�K�.��M��Op�>,E�B���EX&���Mp�����0��g0J�z6��T�y�ף�
��g��s{����(_-��6�`@=-�	��'l<�C��u�ln[뤼T���PAL��Ce&���Lcm�LJS�������N(; ȸ��,�P^j�����T��O��s�1g�dQco�\��;݈��_�2��l�w�YQ&W�(����c�ݮeޔ�u	��"G���q����P�7�%͸
h����ڜ�-��>�^��4�t:1W��ebB3��g�h
G�t��m�'�y_���ǳyMF�|H�\���4�q(s�}�g�>pr@�Y�H%|�L����t�����3L�]G[���RٯKzR�p���:O�ݑ'�M�X�3�Q��`�!V���b�kA6M���C�;J�Ņ!ў��t�����*5���>O��"�^^�^ے���2�tǰC�B����M덐���z�bC�fp?-7�v�6	{ަ����e�ʵHnu�+q��St�,_�ʝ��P7�^�mQ�s�Kbm���J@MR͑����.H|��+��$\�C�[�4Y��AH%�ɂ���IE�S7�P��@A�3+$�WHJ.IgE���F���k]�
r�Ā�	�q����W���V�	�:�%Sx�%9�5�=���Et/��Ӱ�ZS����θO,x�@l�M��z�s2����7�Ĵ�^�ua
s�bx�h��cj�<cn���S��K��^W@�=lq<9��drf�H���.�!�N���/��S��X