-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
03WZPm9FpS9m5iFT/4/jaiY8k86hJ4JfRG0gYAn8qcFNUlOMRrJ4iI7N09CEpoGWXsMfloTi/izL
YJjRYai1pnLbUkGnSxTQCJMrVPgInRWmb6CYTyq0DNpmbefwHDjeXoS2k4korZAJLaNAsiMcpOWR
Xo7gG/VrpCQZPWTZUhbp7dkoDuhHIoZyz7mXLI4CC1IvQ3Fx32vE/TpyTjZuv5x4cTnvpT3e/zyw
NZ4/rWzTUPPKCMXleJ5V84eY8o177ym4QD0ps3D/q4rKszSFefEaxEYlBoNydylb/+yhLOC6xH0L
9MLk2lt0G9cOK/WJA1EK2JWT8dwFnPm55slmAA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 6512)
`protect data_block
QOBwdcmOK/p3Dh394ReHRkjSvq7f1fgdDN4n8yxbRz7LDbr5hz2AiPZEz6kxnr2mX9v2wlpi73ti
tkRt6sFG/WEJywGbeDvJRJGHb084Ige8A0H+X00hM+dvIcOj71ZgOhwnPeu3c06rJRKOwsaqh901
ReywjIHbGjQx1XPBW2qU5uUVPAktGBfrV12KH9Nv6KKrRzeJzdQcUggOmySjiELK61V+nkBavb6P
MbMRx1lOw5S0FzPtRLS3H2qcEa8BQ0Bd8VQRStGNfyPyr3cwsew2CA1QW9f5WgCwLWqllHZn+mmC
Mah5ETFqbcu8LFoF8HzzmNvMMVsajXY7FNfFHfyryt4RdXneIoRuiEHp4F6weKhJRLdJkc5u6qIU
hf6oI3mP3CkG5SLz3rhiOUuI692levjQHDud32NL6GJXESDluUNcoS/2aD/1km5KycMAGP+aIS68
+6T/MrVZe5HoPSOGcd4LmtarVFEupBKLyVvtYf8cqmIJV/FpPB3BCLwMkuYKmxqXAnmcwAdOrXwo
VNVu0Tgm9Ox+HfYbovOIkoauCTQ61pt6+QOoHIF2nkrbko/vCSrq9PZwNFLtbEPEoEAhKp3D/o+C
XlFtrgL/U0TlOJNds5F+xbuZysr/W2I5L43OFNfv/dncbrLLR+eZ2n+GPvQNswfxspL1okx/LUXT
Br+iKVvFDX8Ecvj6GwxTsaj8hvumJRkXsnzSPMVhoLkjbmqVivaOyt7JE/iNDC7xOI8A5HkIbMb6
gp3dAOEcnXP6Sfqm2NMvIw1ieMIWsJXPTlqUyJtNv4kbdCMqFXyjnopI3n9CgKi17Nvs8/gbiTs/
JukPChRGKsAOdT5Be6lSWEYWdHej/KOH65rNiUC+FTH1gYdLfWaZ63VY4gqaakZ/hc3BoTU7iKm4
mes1m6dJlmb5mEhaC7JzwGe2PjY6fPAPTiabq+VdQTh/W/UogDdm15Shqpw3l1iZhb/YX6GlULM0
w7JCZ4MRDv+GgBHC8S5Et3eqmw461irqu8OvyIl2iviKNU2Q1BiSU0zrYsegxTkZ/N3Fm8xTAQbJ
a/PaaIi6aKrnLcRa+TrY6UfCOA2gKEeucFEWDPVNWMXIS22yHreyayDaLJ2Vzt5SqtPbX2BscDkn
eoOABd5hJAGo5CYBl68WIKy4jfBxO7dEnC4gZZg6l+DVBojhL4iG5pJLE4fuir+P2J1C2HpMDCYJ
/+yMV1HtidkIB/FCF63BS4Ob9eF2p3t9B/YVwWh1QLHElvt8nOKMSZsOGsoPPZpL/CDzClqSFGzV
gPFhP6ndo1rrNEiHGS9enH/Tt57BWegsjw1122tvFk/BjoyP1LcoVBmHmRRqLSZTtqypsBmZtUuf
GXPtD/AE8b/eFtSxYORmEc1rIl9ch7RjMpnFRwDXIvFY8vOgPQ92/PKn25RT6NJLnrrnfwJBch2T
5fnLBalwQU1V9YaV5C2pwjyFYH2MzhjBL7Tv7LMF9y3fjn5J+0SVh0Meu7DQtXSwKQVS25gGLovX
1EOKgfXy+mlm5ONfegyv42SJ5eGDMd+LxUq8oNKSEKMPpMFZ1ZQuF+nzNW++o4ui148yuVv9fUWc
CV19TYE2Zp592K3jzc4opmcO6OUkoeWW3gawDCiHpy3FU9HnvNFk1ajlxSNCXP4R0IrvBMbud50/
Rq3+b8tUTQz+FIBPnPANNSBeUS1KPcV5kG5Ehd/BtdvHe996dFSOf2sW9NFfEPOUNZaFS+EomWcZ
/ymv1lVh9x62ZtsOiubD9+SQ5WBL+gPSP1hFVFZx+1Eh3vmr2kurzVFLFPhAOoDuQxp6Y+9I8XKk
kSykuCH3u/4WtN70q7zSyu1NhovDpkbiiks4HwnoRrvMGBRH9BWIEegKBFDA237Jq99r4fC4zoMq
HOK4pEFFcf89G1/rUdCEkI9CC5gVYNZWQYlarc2MRXiZE2XH0IuvG/+ste9ulcybomCl1LO5H+0X
zlF4jfJ+5LD+fZV32ENYprsU3iS1mVVEpnrUpB4L6dazHPcr9B/rGi0J/kqKGe3a23+aYjYexWTp
TrV7dgm72KYt6osWbAnRLGLw7TQzkWxEqO759lxZlgkfHjXhhTHOs96o3wCNbjkTt/tJswdIa/kT
0MisiuP+Mgr5Lvdl9Rw+0lCRn5OvncX0WZC9ttQkdU66xe9JstecTO9AfCKUuksHg8UgbVZSy1ls
lOVCn9tgOyzSF4v5tcXmwSvxesMXFnEfdoCx7SBQKTq3gkVfyc7Ea1UWNJ1geJMvFRSUUO6nME56
IsD/+rHjzDKDjSzXPYS0Y5cMDINDwNoW+L7pEa+X8WFYul0ZdFUEIEKiUqEv9dFNfCaQnDDYjeOJ
wYILIefEFqwfsfb1unYWDZm7WYp3UINHLHMX+MiYouasM3/OfMS90YeFfK01thb8HyPjAXhisjoa
PH3r/ZFE+1Xyu5PQbqTm59Pfsa0Ly49L4EQ503cSeEDIbHNx25ZSo8XP0gPx9/23Sew6e0MeXf7l
iMoF1RhDdjUafDW0qMSOBy/wobSe931bz0FMizdTE/z+Ro3f5a09GnXiVQDKkEfA2CQFoqvE6K2g
4o6zLyqeB027sVdmG4nFVc7zH0XwBItZmqdl6zROLksTOF0lbXBjjbnWv4E9uK1aLYQMB60vnJ+8
H8iW1rAGjOGiHjl7CRIRAjVJuUFq6N82gPvfHlxuUHBco5/XjXKleRWkf3jaOJWsnN9oaMs4J0sD
FLbf8geMMfHxRLymtKp3z1P+9IzpFWMIoscn1Dua2RU4tA5skkb6TIGxWthMBoHCkk+1ivuTbGbA
i5UuDWP9inM/0ZwoEiZ9fWnLbkQhKxO47kk0UQXbzcLe90EU6T0OE9WW3UdLNRJkWoM8ho0WUyzo
ZqUUu4bO+zNOgOcEvfx3l3GgJQlhkOVT6ReZVkntY+cV2zpelq/eBjqaZKFQaiIEfwE1yLIMOsjW
BA+BjlqtP9HiFV13R7IlccvuSj7y7O2RwL0SzGKIH5oRaViBaFk1Av0Nv90SIHZI/H4yZqg8GjU1
JzOcBMEOd27QdVUL1Sqha03uoMfh4W9SDWfNzT2OgWmMji7jZ6rD+zLl/7RdZf0uGDnXO8v/96iF
KD0ONwLVF0Ha3Nj/XZrXn3yxPgGSJ1eii8ixj8Z0UmqhpFRqaOKiJpu8PgQWfzEjvupQNmbJrio3
9n17sVXncFf2pNtT8Jce79ynUxSIRBRvNLeTnlrq2Y1EXadaK0UnYEY6nANqyZVBmzSiOh06G6Z/
r493PsFKe6ZeM3PghrKGEpbDNrHMYT3iKvBgGMpSsP2mHmpamRObrwmTzqStet0Oz+wklsIKoEbI
/YIDZOp/Yze9BcX6W6CiABWGfOKOUafEPq4nbFBzdWL/q2OQi2HT84TosvPXoWWM0DRSAXvNl41M
vOn6+r5C2DvW1sW+okIbUL2HP3Alwuh6niKA8mh35EQWB5qy1wjWkyFi1ciWjAUnsScAq7vGD5tH
d1wRIEz0pudqqIe9pTjCCvPgmXkaNetuRttJwi9hNn7E8yHOfYyBZ39/NeqRtIDr9TacD9Wi23sD
dLVFMau4PJST94H/11mttEdcRzzMMXUlA2xRPwbj5LPMItDcnDeR8eGmWrtCnyxeLIpe5Luy8pxr
BybBQpfQKWV4CySP//NhX/iY03kRyqXyhu4koXRrBGlv6IqTVRuo2ofoenfga+dl4wAd//74co6p
R5UebIu1TT621AAcIqAMwIgR3ObdG2Oyv4MF92zYJESw/So7TQF4c7WeLyhAMbLHb4hiunn2dsFe
DS8vBoNBB+uSIObMaxgGOLCVq4wjJtg995z/45zg21jmTi9w28nY/efUAZvBGZwcscRrLk0+UqXK
MaY8HQc7i15AWzWz1hguDDoM1owOTQQ8MJwCKq/k6qLuurtoQecyx1+kFdnlaciaNrEKo2TVznBS
+QLe5H4V2vJ+NaaaKb5cuUEGWYr8GaN1YLiMFzB+zzL7IDrAsKMCc4kEK7kjjReAad3bOjsqKDyi
h4BVQEuUd5l/XSG66gj2xXAGl1UZ/ZpVv+1JHC6TX4OYrzU62YrLFm6j6/9UhuSZmkQPcQhL7x5r
Z++vBwubVw2TSrXpLnYKFpJSiV8Mx4CSswLfC1ceF/qHh1sdJre0ju8F940KWJXd1hrtyeTopUlW
JCUsbVdW9MODN0p5/G7E3aF3rVSNCg08eh4Lxx69uREQCb8OsP7fnNk9NDq6qmV1YNH7XDgJuLDI
5sFGUAwZPwu4avFn7wPI7ahrJoY0LgRTRljX/exyY8lwSlh+49nHUMlI1KnwgJ0TG+VkCEfLJi4l
Iy/gVM3gES8EPRmEbuuJkC33cWkWe6rQyH+1exi+aW7nhYmVXV5i46DByTOPAsuvoGBMnamGmfX9
fi6EFl8QvAMBrJtcx5dq4vSzQAgsVQihgGg1yURwVkU3fdYOjHIjLOMvv7tWjAHAaiX/xOA4asvV
mp8uyDHwXbarTMo9Mox/o3KB5maW9kDtHYnFrTrS6PfxzDHAmuhP/xZtp1FQSxkzRx56Lec5uRw9
2Osn1crRRdA/7FTnZSadS2Ybfd9W21qZ4hxj3Vg52ZG/J1wtfNAK3671BhyF+GTwO+aDea+MKw4/
ZGEa/wDBGLT6yGNW5+xxXoBesOtIJM7mtwJR0r7SQZ/wFxxXqK0Td4g6dbm0weUNWpHLtAoG131z
3XTOVTsI44rHVO0oCTjkwiKyde4rg1vx/D9mDM8CiKkKVCdJww2c0YbpfmxkQapBGWUoF/C7kcLE
2cJ+42vIwFcmwcLjBGv9lKr0Mk73nxeh6jtjZyUYI55l+Id+jK3TUSzmnrpW1h3R7+l9TW+jQGP9
tUf4nizZ7I7wM09bi2kToS8hOUpucfk9Tpz8Nb+ECPO5J5aNAc8ot5FXsb0d5o3aIBO46AsrW5P5
Lv7y31Jd4zgMVp/pJBDJqzAVPNJB/LALlUti3JbyRWQHsz2hqMlF/W3ovZyFiq7MYJTUMW11CEiQ
OWRtVA4HFj9IsCg/9gFSGbckUr4WJSSEj38yuvOqwSXf813ZBuc9x7F3ZXdMvuqEkVp/dGvctHQ0
dfRMpId8qfwgMXtN02r4mY1+py1qY3qxIK/QuhsOddVP8NNrkLihtcVJlzunSR8Q9yiCFI3JN77E
uTwZUPQEPGUB3xHMoezf4r9xK7xBY1UOjCagNk2+y59KacqAknL4zqShwfHV5iW0A7UvzvBcjmdf
CS44QxmJotc3cOGDH35NWoHMeWHIS0FnB0MN+TygXbryyAqcVi9d+s3+9+CRw7m5mU+kzA65islw
/sik5nKdNfKPmu3nUBzHzFb7JEE2RYMiARCH74/Zkh4YUnMSDSb+kyypv2XuNzE55eHe/a4QWMMR
GVfSAxRTmKB/bnwWlBOYh5gReE4+VOsFwAbngMT1uAlyE24E46yqto8+q/LhCHnmbZx9lkC4zxpG
Wz79ZBmDVlcdgauO9/tdobQzidDBcM3OjiAkDBU7or08KQapHFSC7S1fqdESeQc2veySmA7y5s4u
3oPttG5fTOMzR5GJXU8OHAFm6NR2RhFyKMTzbQZw4MpqDG8CTgFQkd8hr4bpkNf+HslJzBAB/soW
+b/BJODitkJJDxinT2WO1NtiCzA5qWLnILjZvGSlqUkOXyJMmTJo/SxV+XvCPsKaey/5Crew5Th4
rK1XBjKddxyXO2LyLXiDeLW9YRcjemDI/gwLinDG9QH1PPefVebOKmcY90yz8pitmgMwhM1AZgBT
AY2ePqxQeP5oLSadz1QcTSnxJUXCQrC11xWvDTMfg2sYPW6SJQ6y/072RbDBEbYs8qMk69q2PsMP
mqLbgNxY72qBW2cgulTrq0o+yVEu2MCWbyljDFs33TX6vP/UgJ1/aGe7K9y/mZkcUrHy47bMmUkQ
qakHcCPGsN/4PUL0p/RzWWkWF/oTyMyiIgEnfJh/6LLOdcP2BpruDhkTR2lksQ/36moEIKrF1xFv
lmUSbaM6N81xMJvsHAmlZFpsDVphEc+imClKfs28p5jhq49PUQ1nL27y7GhaFxQr4VrdLVtbdeDF
cDHMOmItZ2twpDF06fYd2FWLI1gW/Y8FGKaQ318LQ+y23RKHub865dzVrulWsCtMWo1jFp6eB4Nl
v8o0NL+O4cufe/4CX1UjdZC/+tdHOwYMTVeItaxjAXfjVmRW1pG2vmA1b6wlYVUmTZMunYM7hZlm
ScZyimKnZee+L1KT1A/uh8uSuJYCsHw4jaDYh7YGl+qL++tWarj+4+kWdWSv1CpUjjunK32jMHL0
NqXxtJUACJr3PHalAaYMIt28VU3TKM+7BmRWRO5scZRaELkgVYvcXLvjuQ5Ggc4c1fPu9v8xLCOM
FhKVVmQ0olWb9WwYYWLY+3QlgH4IeU8SB7vA+CBSYHLZG8ku9//+LC7YiVqUxRrMy6ZSza2c16wV
lNhLs387Yaoe7VJOotT5sMjwiQ5MccKadtWmae/vTpYROYP1g4N/DZX7rl29eiNO9FvgiPuZN1PL
XiRuMzSfBocpfec1ZcioLSf9tPW+ATMk5kVoV+SoWG4EmjuGx9pQlALkSFfzgwqBWSCiK0zuw1Z2
duB/8tS+e37k6h0sQDeRw2ESu8I8KKutoegZtP5ZiRpJ923tkanfGwnzQy6Z9cPWfexZFvP9hUje
tCrM5XMLL6dW1TsGMldcpMspvxfhZQQPSY/um7H/89y6xBSGFScrQzHwWRogRiadEKM1qsQ6HvVr
FbegfvBZwP3ltEJrconoN06xCp26uRdCS28w6pItgh/bRgi6AV/kKtT0SGCG6/LpeCGXQOnddcEn
2tkiYnTou5sIzG2EP9FCI0sRNbCNtfwwI1dTD5vCiZ3wdcaRr2sWtBRZSjrQe4I3MOJObEmAeDws
B9e70s+Y7aZrVwu7hhK4FVk8ss3chkQvQAlUfbFaYVWcOTwAreVAvumlF/luvZbmXeDJgEbIzG3N
ksTH4SZhkVnqNvPu5lnEwTNWiiqrDjM9tv94zmORSishZ3vMr4gmxV/7v8xi5lKGuVGe3uJMKHYG
KD4RnQAMA7voPRkabFix5mT15FyGG2SS5LhzL6jQvZIW7+/Xm20EF8JtbuufTy3FrWIhAmEJmjSU
Z2hnh1qBf9/4wFlzCqrfoXFGkvUWOnt9wrGSyPRLIx7LKujjmWsMNz3jZLLrDQkVGIfiqJxmyGRz
7eCqfN4VxobvMmcxVLrLKegivIEXCPG7Vj2VFnFOljNmgWZwC4szo5/gBaL71f1iyu4r+PTS9Oda
BWctwGVgM3dluH4zRIRS5sMp+6IkPwub5ASxYydrZfGOIgXWgoHGygi4M/Xh0aGsdYneAQ6+359c
P1EblSQB/fn+0Nu1iNuRDZJJ2OhowlG4Ct7NC/tHvg2boUT7hK6Ii3o0LswXx0VEWkPOy7BH7UON
2hMaxEvdXylvvXnj6SxuAyh7xKE942CGJSoZWzUajy7mqOmoUgvEk5UR8anGp5y4QUaXX6R9dtZL
wTZ4EoO1fLMVhNCWeVd9vxg/yAuJ/pQkR47CNYpP9FzZyMlKR+LnKam1AqEB+tF8XfxxPRilhtZK
tbLp/fNKj01G4/aV8tQavakmgICFXzmwXmBmikh+DQs9rSap17dayBR6NWAKFqSyCEo9+wLoTejh
Zs28DVJbPQAeGImr/FsUFjLWRfX0Vqf7PlxaNPP3I0BwG8/QRMVnDCT4SeOdKyzp1E7WwRDvkKjL
zkdRWJttcTYfOqGBYBFuQixTqgi26BLVtlsR63NmKw3dlhLYc4a6eGsR5DewTJeQaaFGnKE6TXcU
bKtTjv+CSvIwV+Itp/GKZqp5iwfOyobuncAmdxMj9Ai/ohj6Wvdqer76Y/k5YZa57Dvi+lDX1Jz8
GnIASp1z6L76R0J3J7Ov7laNaKt9BxCFk1zE5W+X+6EgOm88g+sxPT+tmQPf7Cgo2w9m0xURbPXK
Di2krAayEgA0+LjE3l9uivZX4CKy66fNcpmNKaCMOqsh9CdMrsICpNK6FKSAl9S+vjZ3wyCVXVQe
TKR8WsFwwu2zb1NlL/of6Pa1uIiw6a4MOeP5Le67q7Tpllrb7GK36CycmQvD86jx0KjmEnzNgToq
hMdzNCoUAICQtMY1jj8hz06iwXkSqjv3eVFxPpS3BtQ7xca1XA7Xx2hsogzGF/rwN9cAglOzC1xq
V5Aq/13DUwdhl4uamfrW5n5WTA2yjwQMtjE0M1ShqSr3JFoXUxy0r88VAykEFihfkq3ilot9Ea73
SbT/nD2tql0OZ3oBicyBQJy3oTaYRh2v3QpQVfFreXjY3I1qCvINkHkHHt8zKEKd/8B7wC5NpUS/
aO8dJ6MPLXigoIqv2hJlL+7ELYZznTHDZJE224ZsH/3I5foopmdmrKhhwZFWXQN+t+w7I699r5uq
g7f04Dz/tYmg3TebrB0QUypW3qw5CRK+9yHqIzb0Nm5HltFinTpc30I/MkOZs/oySYaMy95Y4+PR
olnL+fLixi3g+jHYKeUNMIdJyiDXOr9Y8vGH7z26uAu+Xr7KdE4xyg2jgM1hNr2Mpl/VSEXaizIM
mrFJ9HSM9S4U07qlAMzdwwX3dSVOYAjg45MIGT+/jNx1MpaZkziuvWI8qIo45r00cTtKs08JruHj
WO+xg7QUi/KRnBQVKg8=
`protect end_protected
