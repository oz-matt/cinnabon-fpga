��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%����B�/�u�'N�jA[�Q���R�����L�-���ZSh�O{"��H���,+�Cp/�3&��1wy̑�s���X��5�&-}�IvDZ��ϡ-� 偙O��QZ��~rL'�x[�i,mׇp���O�I43��4d�,�H�����SN��d���3���r��m���̨T�I;uj2Y� Er�*p�Q$Gm���p�V�`�2^���,hz�<p��l�Bxt�5��s��\yq���#�@W���f:m��T�	,*�񞭋����_��㧋l�	�\�:��uGd��PǷ��N�I��_����Tuv� ���us�(H�~�{2H�:Zor�Q	#%�3ˠ!��iS��95�,?�.���/�F�i{#���Tp5����Ҥ0{%���2vpn���X�����@l����3dc�ק�3	�Ed&3�ZN O���z��s�yxӡt��v*}ԫy nj#��lc��m戭k[��5)�A#�����8�!�]�Z�s�M���t��w�!��'ÒE�rv��Ϝ�c@<U��\tq+��&|�&X1)C�����r�A~��B�&�����s�:n{p��͠R�X⺂L^��R����c���f��J^?��ܣR�O 1�rV���:��T�4���AD����˩�F�w��)Dm�O�b,�a���1$��c��7t[i2>�ޔ0,S���󧇳Ϟ�ᒨ�-��}�!6��Jyv�醊�^_�(�H�(y^����o#����X��3-�k\8�M�T�"`R�DF6ȕ� �,5�;Ҭ C�k���1\������k�t־9�}���� ���QHF��"��t�9 ?��{E_�7��!����]H���L���V�gјmd�FlЍQ<aD����f�x��N�6�۠��Km��,�+�Dm������Cq�������};��,���cb��	c�K[{�j������2^�d[3�k�t;�4��wߝ�s a���]�#3���Q6G�*;@�@�WX�����+j��3�$�K�B�V9�q�{�0�J��C.����c7-���7]��=�HLD&�J=G&o�rq$�
��>X��࿬��˹��յD%��ٯ>����{V����N����Nr+�B��o�}�g`�a(<d�t})�(�<g��&i���~Al�-�vq2�}m����c�hj���k���x���NY|+d�?�v���O�W���p�D��c��[�<�~��j�1����>t(����N�Ꞝ�I����mÃf(��B� -N�9����l�%F���0Z�УWAR?����aNƃ�՝]C	�׀�����V@r�u�/х+�JC�q�K`���S����	dF��y��v�+�*�)%Ck%本�����aȾnO��55�e�5�C{��/x>>a�%���L��G$�
��n����h���~bx�{}7�I��(�C�ӵ��}K40J�[m!���?����Ĩ�(��5�Tb���Yf�텲h9I;��,d����W.�y�uR�D²~��bG��H$��r����(�S�f�݆a���V��h��mLP����>>,6"�B
ȁZP���I�kT�
V�e��W83��'�O�!�h���]��Lۦ�9D}����_R��C���R�.�4�w^���m���!����^�X
�82� �e`�X�!���l�~Z�����x:�y<��t��㸡Dp鹏�ˈ�<��󅟇�E�����O�wW�Z�]t�\	�4���
���,hvG=�4fGB��,��fg���ڄ�U�A+�r�`�R,��%3�+*�����5������6����ޙ[P���a�ʊ4FP�_���J�NbV�S�Dn�CE%/b0���Y ��0]׆���L3�٘E*2yx w�V<q�jnWF/`�rI�
^���<��娲.:&si���YD�M6�A�ti�����l��۫�{_܌Pt���FH��(�=ύ4�;���+��t9�/rԡ�5:�NJ)V��^-?@���<	�M:���|8c���v��?�3�am+�����,���q��4V'��=��ю`���SkN:���zmc!��P��\�\��:(zm�B3?�,}�����Ev���< *^���]X���v�XX��b�P8S=��Ε�fjrܽ����:��{kP����OF��{;��Qr��gWKa�Nu�K�<���GR����e�� 03nI����4UP�~�ŉ�B�mս���	#�'hj���MCR�!ّa����w����D���45��W�.��B�*�}�����qN��׊���u}_�3تqX=kV<��-��d�#t���q� �v莩�d[�i����
���"��=<8��R�F��zr���/���L\�W|@��Oya��*�\���Ŷ�L���M�*���}�xU�1�=��;���[�����g֞a�B�;.�?ui��y�o�E_<k�����#6��a���V�y$)8�u3����A�O��L�.�}]S���(R$�+վ1���
�͚��\L�]�X6o+�lj6B�Z�.��XX/�/O1&X���6��#�6�UԐ�bϳ9/��ۣQD�� s���/�@;h�֐+���4)/��z8�F�b�?�M�X[��bZ�jyO�T�A'��3ٽ�G�?^��3�u�\ik_&,��:.vΑ��A��b ���B�� TL_;�s``^��\�ڵ�S=���CE.c�����Xԯ0�ݸC������Ϻ]syZ���3ĺi�&2C���>2X-
����ɋ6L�
�^�(��dx��l[�/�k8���|�wȓb�3ڠ]��Tˎ$4o��ͫ(�2*��r�7��M��$�J�܎HF6���6��o��zP��-/(�k��y��b��)U��쎦$n�<@�Qp���
���)x�rw��.W�5B� b~�&;d�VL�C߯����te��Y��6 W����h�Wi0ܝ���
��� �Խ��G.�h%ҍ��/��tee)p('@T�W�_3���4����K�8k�Vem�ĭ\�_�'�k�)(���CN��ӾCg��C�N��@2AR��n� Ѧ���W��Ȫ�K<�/��YP=�*��x�:�.����T�4��?�O�jr�w����	���)|l�5da��|��i����rvDfӃ>o��0��:u��#4��Q����1�Y���(׷0qLa$Ynt�}���:ug�יG�0}=9�S���������V���L��k�jk�}�1Y�m�)�H�]��5�S��~yw�>��v5{�Q��C���Z�t`�>���T��P��� �OL��=����e���'��*�'��},�ħTēg;Y 5Ǫ�֝3�(5�H���c�Y��,T�={���4^Ia���~Um���,&ݕf&�ʭ8� �]`'�<��^F�d�_���\"NF�*��g뀧�3����!Y@b򍆛��Z(����v��t��K3��������<9H��^�!a/�����p�T[K�S�L�
��N�E�P��-����������l15[0���IxĲP(��|BI,����� K�P��˲DH�a�Xe�&��<����x�&�xh����3z��Ml,_^�F�z�+ym�x�3Rr�m��d��΍�S�e�'п]㈷���!�*�����D t�z5y2�;���dO��UI���U��H�J�������� o�q%92ces�}=T4��F:�H��X����\��0�x�NYJD�U(�$�۳�Z���!)��"���e\/��r*G? �##δ�����*�d�
Fc�s+O�h����s������_����cKdݕ�Ҵз�YUK�b^i���⺖���c"�UW�RG0�$>���`Y�Z�{{�jB��F��T��ZGw�N����X�f�C�z�z�Ӻhe�S�X�zr|��uX8K�m,��⹀�_ѕ'`8c�<�#���z�������%��닡�?	�o���8����#V���bl����Rӟ��/����;QT��X���IY��7y��ݧ3��� �*�gcp2�*kd���P
��g��� 9�|0o.c�Vָҧ��\D��v��(��*k�V��@��K�w�AГT�uyw��>M�te�|޹:u�>MA�Fu����A�i>r0�=����s֟|��M��p�ܲ*8<�3�^�A;�l~_���C�����x*�A@PT�5��4NV1��C"L��Z�����9�[_�~�9��`�y=�6�N�qF���造Td�$R���B��j��7|Ϡ\!ڷ'��-��c'_�;,�21;�N*d�r2	 CJ��|��b�T�3Q��˾��,��q	��;���?AI�|��U�)�[~�Z��Yٶ�h�פQ\*���O�|�Y�Nڤ�|?�z6]V>��nj����G�j�P���d���cD���W�L�'��ucvu�y1�%���7�]���*e�����-U��)���N'8`�`zv��z��u���x�-�w�}�%��30�=l	H����@��;`�*IgS+*Eפ�'KhT��#��ȼ�PS�N��K&����$(s���h�;�����Mi�y3���@Ґl�P�0;gi�>D��{�k�խ&(B?�a���VY�\�����&n78;��L"R��]�eTdh�Iv�����JS��J�� u,�<��B]�=rouƭGv>�b�A0R�t��K�`�qx������� ��� YhUG
���Uܔ)�ќA'��vV?6b�-�}Ћ���XΌ_\�)��|^V���R�ƈ��vxO��\�����ۯ���Ix)[��ld�Dȝ[�F�@5���"?���t�1��?�O��1_���F^�����b:�`-)�p��o��F3�X�H/�Y����Ns*��˫Q7�$�
���b�5��hc�?W�����Y����p04��4H��6�A��� u�.m�m���qx�
�Sn'z�kK�Oi��xu�oP����Aw7V�;/a�E�����4�r�X��{�i����m�y`��8�z��nQ,�M�Z!����d���J�~���3�4��G�{f|�dc]*�L{-Ť:t3��S�y���'{2m�J\I��S?1��d�.�P��������t�h�ff�G<{j�<'�a�\�{���r���,[k*�-:?���ϕ1o���h'�����9�z�<Tv9�/3