-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
GCijy+1L7MVWF4dfqQHLCHHk/4LhQ57QhG9Vd5LwDMl/8eA+BxxUBN8aVIwcc8gxdL/ZbmL6zGb3
+klUiN3AnwEDoOHRgUnWlHdPeVozI7c+7ZZeFakTionS6Snp1IaQGE2tDMQ7U0bgx4zwaVNevryY
zog3ryA21tM/XZRw+Z7S3sp4P7D70yoFfXfdVZkDGl0XmbH5SfWIaWd6vPPz2YxcfB5JXH6gXafu
L/7m3ZGluqAxkp/jaKAWAE96yzlaDcR49AAqLUuJkyqE1Pqnx2WEpAa7xfxU6UnfLn6LD5xVXiyr
yeo9vzfzZA+g1eWRgLDtebR4J0B3MmonucKLJg==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 25280)
`protect data_block
7UTfQt/EMqOQi7Q5cW7rpxXqXH8h1AM8a+00GDcuQWRhzEiRmGWJhiRKucNJeqJx8EiXbBtsP4Xk
V5uWd9ir32P02svmLQKdhaUjzF4L1UgVkOWurkC7bd+Yqr4I6AG+R5Srx8rmIDcVPQg6gglk3RHy
wtrGbzIoUZrIiC+JTPBmcccnpPKW3eX/aXIMpjxp33tfXYARHwijyNQT7RsPu/sAcayFqAg2ZkZ2
mpoJBIjpfFEJ/zoE2oxd95s0nGGbqDfvAQrmvRTG2vNiKt/UGVfeo7qJSuhK7f0ELOazbPX+rKgI
/QXEs4MAhEZ8KMoGMApoAWIO14Pk7C671IEOld1ggWuFRgTBtbNnYNr3fyfZgqNegSAJumgbgUiO
RDUanGo0wqrYC5xghJaqFSF+5sHmnviHVn8j7n/CXr1VPYLIDL/K57pfxMvRcyzIUUcVtqZ+PlUb
j4aA7YXoIclmUT+IMwJ7LGAUPVsoPcrSwBmETPmElejwLs3L8kR56vA/CfNkihcYuZDEHQtKp+le
6D5Izfo98ILcyAYFd82lQ/G3+FgGvT/u2cZOYhB98Gz9K/OpPbSW1bgw2S+sHTH5hfr3GbAtASCB
WTjT/J9NRtCyyj25qQeQOM3xxYENo9NSQ0tS6qRdKZmVFpdQWwaxkTLQL222oAtzxgm3gYPzFz8s
fAzm+fCAxhe70Ev2voFCfGiWM5LbA9lEOR+QuSROQalttanCxMvZ/NseF34XNVYOWHkMta3ffbNM
hprbSt8MmrnWYKUVY4JcekOgPpA2Av06ylc0yIlIOSjYxWFmzt+82ZFJs23J3t+bVYvUT4IijCXt
fh+NKu8eQg1awfA6NmR5SW9PO2UedIAoswQxKk1z3IK1XAmLCCVzDtSVUwEzCbGP7JNQxMP3hCFU
AHh4+qQy/GcHr6wR1Xik9qJDjALiBGpRDkpjPQlp2ewWSh/L1tHej7WQ+8k84LQnmmybYiyZlAPA
cIdqdXY2xPXB6Rk9dn+daDcLLSQX7mFwkI0HZCmuJEoJNFzLqrGJ68ltR5avpChV/Dbp4lh1N9R1
Pk9D7Lf/uC3v1wgFbpOFZLMpFEDuyaCNZODm60BIt/hlwM/sw2bw/au6Z6YsRKNO623Zopx/IjtJ
ctpYJsWY5TBPNRZZwuqzX4Vml/cOaXt9D1Y9zoHzS5tmIWf758jHh1ST72PiwsO3ss9bq6cqigpd
kgGH/QHfdZ7q/j2neb8AwPNKxid4gyT64yIeaGiQaT6L4rkf1IRhg0yHUE8m1yMCwAiiSM8EXh9D
fZSHFa4MBWeVHfZaIoYIpkcevabKJ+V9kbK6UnosiMIEZy8tz5tcejvg8rpvZVgtELzsgXTRC7kY
TLotzYtJoPfX0hCUrj14fVY+YzsIOm38kV3sNxvZxfTdqxVMknDksZiy51orbfFLUPhvVwvzdeQs
hZKbU/ge0klbEBBie5qngCKL7vU6yYZzmbcLhF2X1PT9YNsH6CzEZOPU5/iG6DqazHpwPQ6Qqd+v
yJHc8RDuTBJC/n8XuygUbT/+ECWnoPVj7jugwnutZxsjFuFHwclBVfVZ4tbA5EMMqGbVP7AL3yTP
ua2YJpr9NFPWeNIv+ElLAWw8x/AWSY4AH7e6RGH3ugzx28ATzLtIXJz7o/cywG7a4mT8LsX3Ibt8
FR1wcWq2y+tOyPpGZ7GEwqy3LUu3NE0qtm2v/hBHq2YcoZOXlHWb/CsMPUEbZSWR8RvqX3OV5ENR
xIekvI3QKTaLlCxFg3TvHYpUcfroXVS4cQ5rXGnB4V5uIAMXj4xHcjjCEd5KAmG9du+SuUeQTako
aUZYT6N4WL+G8EhGYBD/ZH9+uIx9r5Er/+8c5/eTkoo/vnOeJjWFEsEa30Sjr0pvq2A/6Y341oEm
oDlqM2Dr18WMzmIEsNOyehKW4FNDB1zVCM/hL+QydqtTzMpGLVoRH88UxKOdNx3SDF4qY1Lq+FR3
dyK4Zl6HC89vp7ap/pbsah0mYwcaCcbdficxhR5o4ZDdtqFSgP91GeWrOWPkJkXmioLBZe6QLi7s
0x3JlyvfppY8jDkPQ4S2I+EtLfWLWTC7VyADCk4MtdtZKRERAo7G5lQhzKEvOz43Sdn/AL3KqBIN
0aoVBrcGKsZd/7h75B/AJSPNdtqS4cyOvzIXI5yrCI+Ajw3ZZYn4FB3Frls4OeUun4CkzF8Rivy7
sTtKElAs320pqCEyB05Avj52exsq1rA+BeIzOuY2cd2VAqOW9Dl+7dEaRnpXR1jwgjdf7agqeng2
J61Y/3DjcmsOmswjDO3M9uWNtSk9YAKaWyfzN0GmbsvUJv0CypgH8txqhRXPbv+auaLo1xFZFCKO
eaGE3wRyo4p6QND5ouZ8tQ8yrRELezf0SBoTy+b/eGvOa6qA3akJC84pm6DQJ2ZyKFZYWfnbF2CP
Go3830MweSLnl/f4q5JJgoQEH4hNiC0RIZ8kgN4YQNdFuVgFArkkvc+cQTFNRTqYuIUfYvXMLOBC
GlE1gR0kmFAG8h/eF1iNGhsWoSgnSdtsOciL7AArsFrjdqgiNDe3fc2jILTuIPNWwyS6O/P7VvhS
NfGa0517LCLZuH3eVPb4ik1tzuwbTlt689AxjziPmA8psQ5a99tFJ+49Kd/YyFp8YvMOBW0KM7lo
AjUbN9xAERnHtVBQri40vH16XvXj+M+tfHAFZx+ZVgiRgt0pd6ltVCiFr5pHXgYQLLxAPF2WoaBb
uaquDJ9bCSvm2nCKVSTCbBkGR5716RsUvIBtrCE3Mk/fCR3DCPheAUVGbjoLS/47rHVkSNMalNil
pPHsD0S9uHOPTZ7ifd98oGOoFu5exJdwGaxhCoOz1o1L3zwLMrk26mNNymXPzfLVc4G/My/r2l1v
QfbT118nxXp8yWw+lJKoDzt9NwSGOrtEvAuhVAPwEgEprFbkATZ5C5doGZxnrItqAgdNGsNdbVES
ekQf3fsd7nRSKyb6f9Bhcl9UWLszT5io4i0V+0//2LkJ+IBgIUqzG5qU2WxEPMS9J/KFB2kMGGxB
EAaQ4RzOgG0ySSGooYBGGNGtWL7rWXl30Ia3/Z7BWTieRkqPvsGvVCjEerfad9ZC+0JmpxTy/AaU
ZzxcQkzYrUy+NWJOnzEZ+LCOiwwI1D17qNY/bUe77cVbD3fnMT6O4/tszl1KVSqC+s2LK6bouMUh
zkQYmScu3ajAhlrP+epuPpd5VQiSJZ2F8AaWBqKGElsC1wsy7QA4n0Az1O/Bs21O256fdgl2ndYF
IvPcSqzgd9T4DBqPw/sl+hpOjbag8H0ayuuBClyG2Nrrs1DAJYVCNQnAsf+mwf1fe7lZCgN9b0Ku
A9L9U8l7PUdvKelY+rfwKl53pWCYQb2MzWIqcGxuK7fVVdrtkmGvvoEVu+Zsnpii8YFTbljlyKjX
F1vgYAd+jInh/wSxQT+fcKasROkiM98dD32VLJ1KcE2ks31DaApTpu69xtG9GcpxH116J0v4wZFP
4zpzt+axr9snGsTHpJH7yi6gwZ4UiSQLZTYSG2O8jv75kqNmAukpB9E/JMycmCBqu8SJHjn4hqX7
U+B5pivHGx9HYUt/kOQ4vMfibD2Drjf2jlZRncgYuzRdvHxeSVbnKf7jpk4CB9aEMduycdArMXnK
IGkCVVSlnYeYwKORIs4QuVSgIBdNibJ0GF+h16ClhxcGc3XbJ1SijZzRjINaEnlcc6XwyyCo6Pkl
l8bHA86GKG0R6XSk0WiqGcQyjerQhBvOEcVsMNkNvEQWDMdhlS6RlrsOW7WXXEmvfqvhogSFP0m7
rhtEWQU590sNZ6RQuvgaS7sk0fmjEB0sB20KlKQ52z2wNmeO7K8DbxTMecLRk0qYDaXDNH8UuLno
h1/h5eJ50keNx1pR4xvI23up4y05uErx8xdJWyW0cIJVtWVKAIO4YdzXTqO8ktIWfFfhjCDapCxG
VJug62Y94fEUWa8xZ98KU7u2t4U8DuriSxDuJYUUIFmcNdgohgo1PSKulmIwEXTAMeS4gwzzmLE3
6YaOQ3NNuISZ7JBoN2Xrawli6ycDFtleEBfxmj9lhn34k5aJV7ppg5fnqjinR7W0q8r/qpYRKdoL
K0+qcWlhpR2sPxe5vJKHiRbs1kWCO0efCgTXbezjJTmdX1SfUAyYu7rFPTvDRNe4bBC808nwv2Wl
+GY45gB65LmZtOhlKYQjN9sb1CGvUHm8uJuCQ3bWzcC/+jNEDSs4+AXPwzdDenjvPVBmhEgipFkS
GqpB2vxUWEfqp0NVUuOEOXQ55dh8YlP/oWr85/NeMdV2vnucmwn7zyDw529PCJ6OfUklbzqojkha
ZgOgLmDTFQCXTvgj8RYkjcNOPfeTUFIvKIfUiQX2s/FU/zmeU0seTEhkeHSZ/e4EFwc6V/Qm0oS9
7gKBHrFvbaC45Adtvoy8KILEh6HcOqjxVcTU6B8QbXAAwbUyKAXgcpBPvdDjSg8mCd7ukJxlgMV5
DUT0IyBZkoEIIERa1fiH9VYZuKn+9sHVybcAr7RvSobPa7YLVuA3KJlPvRfYoGlSSuZl82nHCv6M
kruHq2QBemGJrW6YiBaP0EAs4doNEO+rIkfAejm5W13aYIUea+KNkXkyj90Fts1K1/yTxjTTU+mh
blnvdVE3QNMxrOiH3ER2vd+aZw0Ks5XqOrjLGOFL0a2KIHKuu59ioTotetDLC+ynaYsMTFwFgvDM
61TH5CWAQDX3wSFHPKXeve7bmLgj2TcoSIruyv5YvcVBp0cjHYzgZoFWHoeWDxB/rRbwJkdtVGo6
OUw9jBiTbsAZSIaHBMTEZOJBVLU1uaIbAHuP9Xfbdiaft3x2iA6gi5P+EsjQ+gUhFumeisMatDyg
J2eXyuFEiN5oAnk9xd5JVitj4mZMJA0rbwXUzCSX3BgPU4Kr+7h7fJJqR38EhuaqsH1u+m7kAlEg
L6/8aEPD6KkxNbLVmSPT8PoKpJz0CSt0cHBeBHJUTISOsCJwBC3b3i3MZ2V4z6UAU2OANnenvi5F
W2sdLwYQmZy7RcLBEeGUyL+Wlu7tyL7ZLvIkM8PuMC09wZc2KQwj2fIEAZWYtbHIbElvzECBhMOH
xGmpjUymeaVTN3XjTErgu5o/PkAeo6oorWwq0tpSRch+EFX638oZSCpaKBYU57Rlol2hsTvj/BCV
I3QSDFLz5tXniFjaUdY9TEMaNIeaeon3Fd9/HsPbRm3kcho/a4c2NDEZpuWZ/wD0IVksQJoUMxTg
R2pH0El+p9Qq710RRLM6RLHZUyFlvCboyghTRl+0DosqJF5gSjPGzsxI8TV4z7Tha0PQXSu5YVlr
+GcAR6ywUUG0y0MN3hujNgJzBPhGI7q/US7VDmO9zOE0dSMXeOlAk4qfjhyyLDmgWuWdiFkIclwF
WMWZJwWhNnlgEYDus0OfffrxDyFncRVWOeNfN1XuokroovKDF8Q1JhOAYR8++DpSnI+GfK1xiDQ5
Ig7NA+0ESN5zDnDWn22IpIeX+Ungpqk4wsETNkR5vXfCkH9o5JiAqMCh6u1zV0jbdr1WQM69KNdv
Nh8miZca7Uinyu9o57Rg07T/z43wFKry6evBQOh+fZnV36MarZeGCSIOSg6xWhVhxO25wPxIzVzv
OrsQmu/YKC8fDeMP4NWacQmhCTBCOrBDTYpyNvhbWUIBHxi8ee42J5NlQ4UggeubJK0xBNcBtGhz
tZsIRfGKfNe2Qe24uDv5SwAZeADEVzdIc4/GOcc+6u6lquySVOZA7SjQinj4e1T4nf1IZTzVnTr9
MFHqPQu0wl89zjjJj7jbND6y0kS9fNY5ZI0fXAoOPFoj6BsiXEwRZ5inNnz2W0Z7dGCv1eCpMdbc
czV7fDhCF9Rq1+wP9rUTx7nnitiq58D3CxpMgW2w9nfU9wej82f+gzI02P3oOLAMmCNHt2oTfJOn
mYW3YCd9mi/pHgfyK3Mg2QhaChcGQtAH6ZsU3aYR/F+RVFdTFql9q2IBv+xIpRd49ZMR/4yjp4f8
fnlYmZ0RY3LeB6p4SGn/L8aNk6O/yTuZcw87OP5wsZEeie8NcnDGXlg0ApoGyIUHwS2ILPZc5BTg
JOLwT1yhLEzaWmwBTmETAhMyk5ANyPAYQOt3P5dChqNfz6So4j8xbdXr8HyUOYUAjGCx6+wi3HtK
wITjZYemY7y9asgdZrVcVIoIUuMilOw6gqef+LQMGKWoTrLKXGOEImojJBrvCm2eqQc5ilgk83N0
pSVRloae6J1NiwQwdIdEeAYYipjMBHkVUdD91iu/LHx4MkezO3JsN87CgrHV795V9p7dChWietL8
y72qdNUMGRanxEnCI0DlaILX9/G86GDWTH/HpBBBW0GaNoD6fJvnjuQcPABZDKCzZbk3CAQGtV4o
9UemKxZjZCVOL7EeWuVEZvG/FZ2w75FmG+RZ1MGXVMe7N1Eh+Fha87Zr9GBpz3baJ8inResWZVLg
70/iyMWY/BcNzV/eSMVUej7Id2/DnCbQS86vdaYDgnaq4rmrDK3TbWTPXZb74aE5PiorgCHVBhMA
j3CxwKwaksTs0bLQZd8+qbt2wqf+kuLB4dmq156sRZM+DOLuYn0pEEYWA2NT8BuGnsV2Pmxb4huh
0n3QRFpyPORv0hc/7nAZSE9AndOrs36OnfluOwIKprBjqgJKUNM5M0Fuf/4oGtb+W51erwZqR3hQ
+R/sAYLsxaYSSF4T3vegxB2CzzNbE+EUUnoIt2tXHPSbLUwSkZg7/WlZo/ytloUQC3+0XruBqAvu
/HYcGZ6HNw4/40lDAww7ikyW4bGs901bP6/ZPtH0PbBEldnlh116uZlM4VWQDpFWzC/Hr+BCIBDw
JC4H0kDEeycUbNveUQ/kzpEyLszW83drQnaQheW6IkEfgpUDX44BKdLGkxKvJk+8mz+my9rMfzfo
2kMbqh6oEXohcvEoF83dWlFz7gdI1vcLp9SiFLnIqDwkSRCE+TO6y8sM9jQVvslOPN4TCo86cQik
p1UjIGLh8ExeRxljHc60F3H3X8EdPqevQC/J/utSVJ+PGKvZWWpXOMtA7oYUlF6JjWfmBCpvqQtN
G8MVrctLYbPTEpAkXvkxRwLUV7jrqcdDp75MX7TyKfEKMo6xb0CT2wUMwaApcAJv+oJc/v7Pmcom
PJsIqkizWW3naBlug6yUG4YkoU3+2+OpPCtjFNjovezY8W9aio6XtlKDtpmd7b+efiycsGbGK2bt
4o3qBoDNwTvnvaOTFCrx42G5quvkDkrr8Wl2SyKb7VJiF1F+y5ETRfU9SBxa3gsWK1/m2Aj6EPl7
ZYM8wWktZ9uP5oHTHUnQC/cKRMtl4Xnjl7A6bmCGl2uO6r2SYvBp2PEAyHPYncwVN2socFgxZ2PI
KjA92ccs5DhgOVMDwGeuTgOjAx5gXep7A0HFAhDmgyMXdEnVVoHqpLwQnguc3Lma8/zxPPopZ5Sw
1YGmkBtat+PerkOxFjDjhOiKRWoWzzCFNxNL0KTfUu8nQ0VJyxlutX4OzedmP7Jjw1eenWQmjjZH
NXIAAkk8cb2zEaGX/PSIJ51MQDHEdRCsfKDFW8vZlZbzlYidB3oFzFozL3fCQKGKDf/XCrZkwTSh
SXfzolkBBr8VwE9y1xV8Y36WxgaHFONiSYG1Q5+WYOLOgl1MO5gN4A22UY6Hflew+yZJPfGj9PJm
RVfWBn+OYtbzXhbMlTuHNtXS9WfCFOPY67OfhzxQiH4kK1V/vzuE0FBSWp5TVPwOvwV/+jtowq+x
IbrWKgJIQvyjVF9R60qKUIprT1BWTYcX4SMV6EqZUO3VMAypeOXk67MBF6qNQ25kNP0q8QH7zvjA
8UBSxauUNuNzW5r5Nwon1mUK0sLHZxrlbYzj5HyTPv+3v8I5zRfEsTWQnhBCLSkBBq3rQPL/N8TH
cA/T9aL2sszXdTzSFE8jRrl+wbygSMK97VbMhlJyKcYuf6nhjFH7tLnSNp1WDFeMfq4StYwUKvfR
mcnUSo9PUiB6nj2yBZCs476NnySrjcc4J2eQcr94qBMJpaJmcNzebdI6ZIWDGy6glWudkIvdoRdQ
jq55pUU8xGss+yAnrv98X0pKg6MGbbz9mknJO1kjW1zTsw4IETQ1jeZ5iNE6/eHd0p1c5iaDnXpa
zcB/Xn2kgSFLrqCSBFgy4soEr2JNF3oGducEoT3KJ4ORfKAWVvTmTr9Yb4HFI7WH+w/B/bIaN2i+
9lQhGNKhvWPYVxqB6F7WSrUaUkC9hwZkvmGfwRTtUyvXDlctVqYmMnpBjJlR6cRsh99S7ACJLDIT
/bZMQ6YEaII5/abBteN2+sxUxdmYNW0e2YE0/uSb40EqilJKSBQ3nOQucyQ/6m317YPdGQFJEtzx
IQKwIoJLpy4J0eXKW5cPFBzHVirH3G4URyF6OibWLCGOlaOp0iNhtchD32R4o3IgjhUUD3YBWOel
UL/FwGL6r5oWGFPwfKaqVX3xN0EWpaOAUEoalpES2vtzYB3am3Io3gv0lMZ4SGDyBkkBmUN1gdYY
GaFGW2v+RQnnYClLS1m52kc96K3PKuXzTgt02HyvcgoVdAM2xsTT+kIsNyzpbaYry6VpknjiZ2IC
1okvgKLM9/TunAk7z1RxAKrIjjh1+aP83cACE1T+D1xdJ7MjvrgKRKJKz65vrvdhQOJTOmsj8BqC
WiLXWoJxjfRGEe+KgjhgHckO04IpsALJljXrusm+0mOGl9RMCRo31MWGmEahjlf3yDz9xaV17kgl
PxdlS11B8GNgZMwENRv3AbavDMyxzq8Er8J8JLHpV2dmO/Megl61d1xUJj27xMua/sTj7uTi9Adc
wtdelH7k8Q9btz93WwDUFThvX37QKbAHu1YL/MRNb0tbfp1iVA8uf6VcaCrThnTcNkQDAafGHdVh
tO201RuOGuBFUXt1oghan7HoLFcxwYHOU1B0qpiaYhenxO5Z2kA1Q0Elq1kSPKIg9oIbWGAgJZ3T
8xCqoLMcaZiey/scDxtgJdi07rAjEm/S36VXFgkI0ociz7G9RP+CatqQokZqUl/E7suzw/8baTgF
TMdYrU6ltdd2TpQFRb033caJXna5NoK3nPMEBweZ0dBTUZ6r9hVI0gSfq284IB1QgMQTStTgjRdm
y/x11C9/Y5XNe5BD6mfV9KrWYhfChcSB3sCVvamaSCBEt5Ot2RwCBuP2AiMJOErScCmXBC2U4rUm
aP3F9m8/YmFdHPsMMjA1lyWMPtCDDQyOvMDqKxn0rOSTz4uXfN+5ZsmECCYgbSi7ajdtlWqRzswj
SBWcw3fk5EBwbPcKu7UFTg1M30umf2XHYeh7Rz5KhiL3p74DW/LUIkVsJlSkFCqO18uQueMTlKXG
qupdPTuHxOTEKIxapWYWl5ggJ8okPl3Qi6+Tzas+Nfy+oYyx6SoxnrlBgghIrP19l3neJ2XKGltf
hmu5z7+T6VpK4G43eAz36gfU89Irs5OzcVf4VtxdAp7VpHUIUED7Auyrz5017im3Auhxqiigk+Ef
zfHWoYGRqE/B6orv0hpYsAfNwEbcQBUcek5PtWyvG5JJ/7KuI5XV3b1dYJnZEYgUpaUNYRFf9I+d
v483WcJRXkQUy1/4XSYQA7hfOkkzQQS+q2vKXwLtngTccAG4OeSN+BaPU9JemITTfIiKAYxdeT4y
hkPaFeFgURBs1X7MZBoqZLEiQpBR6kN37J45DKRCK5NHRml3xo/kMkyhdYTjijNhNELKvfRHtyzs
jqxz3Msbu0qyaqoRDmOTh8LTafwjztLMnWyt+MOPdZEe7Ox8sxOVL/BtgeXRWRC/TzGrq/ZVxJse
l1FyHXVzrZ7ESIRKRUsBg1UJGGLWMmtOOKo5v/uFISLVwIqqTA/riuMXkNsk1Kj9iTKuBlY/yGGi
aoXcQBQHbYvMomwmt4GhDZ12R2sjHx+uZwboVw24DQ41YXpyjy3TppC6lMn3DMGUjS4LMrzwLsTM
q35gc0nc6JmnRhPUcCFz93y+w7j9jj+q2+WIPwAm2ZUmzZd7veNJ1TFX44CCSs0EcYY60DLrD5z1
oZ1x0lLd6K1mrnA/JmbENRsTC8P6urdXEZe99jf8KPI1S2s5GNJdNhquRhWL/XbZLxFiWQ6Dg/I2
UjOB3G/pWnnGYXbfCoDJDXmg2X23V7y9fUf7Dzp3IwnUvjAQL1BUWWF1Y4c3THs2i/zle4Ey/ys5
DSswlk/3bq1haq1lxjRif/SQvscNMp/OezUYWBAslLeOIiw0LyfBv7143JH8hqUH3N3feMtsv3x8
wPz29+35PbPKM01eumxOA5Xl3GYImoHEeHwNAVSBHgZ7Eca7ZCuOj2jzlCw0g/8yUxR2ThwVd8/h
vHQoy5f7QsGq9pZ4WaBTGQWHMZx9OiBFTgAvUPISMKSjbKj+F0lP3Az3kN2xwSm2RfgNV9bzwcUJ
7yyB9Z0uMDpbooZybYZ0zFwkeNsZoc85PeyFXe4FAyzL7fpMN1aMHOZ2Xw+A9wdHXWU+bZkHmPep
sIwVw5Xjv7mvIRr0rOQ+G0bk9/t1OK5xBmEJ5f4Q/I03MqTrGIDXEzo4mAT5diDRr0KdmsGrjUju
044QSvHCT0abWIxhXMAbAdgiOs6qsXoWWL55S7+JBF/TxubqXKyzsRVxFHfA3syKIWU0y0claPH1
4G2r+p8qeznjwoyPUcarOLOm9CIGzJI7Yq+0bJPSdq8tMtGRwxtJVbf/yXlIcyCSHAOBO5S6Nl7S
MrHbBxRDRkR9XznodYAyunwv75ef6qXYndYyDDb+goDe/XiMdMoyfuho53ybp0kmna4fTDVZA/k8
XV69ahtFvU3stPQhBDAGlbfmUFiWrhUzlFCRCAZ62o/DeRypuqHwMhDhGIs4SsZ8hm9wdR6OYyja
r/O/YZUi47/kqyOs1jhNjWsMpCpqEpcRZfSVrU+fOw2NbckHrsW89lskdAz6Do/LuvkbKvuqXx1m
Ifmd1A2GwGGGHQ3+Kvo0dkrErxzNoq3fmi6aWS1Fg40YIvDSSpV8iTyq55XtIuTm705ys3J9tX7C
PREzYoMt7rIPVuZE9BiYiMutN9Fi3tX1T1boIkwyRW6vkfi9KRlfWt6JP1x13bGyzVNd8WGEFtKH
+dHw58KpvOU5EH58mcRkys2LnsXAbxr8D4H+JhoXthdT7TGBlII9ilM+atKR15nLHpz1/d0SNTlM
OoELiZmeDYZEogAFD2B0Zc4B9cTnUxzy9iUNT7g/SDY1awA5ILBelezlh+UDcWhIvj445uSIyfXb
VCoQpq4vbRKW+pyathddxrpNsWB+fvZ3CQgLzUuiJp7CVBdnXt/2W6obLYTA2m0aTEl9kFd9lefn
QX5MR4y+K8fCziZh3kAOZxErbqlqM8MdArf5wG8MTmRuBGCSajNVo3hoteD+qiVv/QdIymsIJqKA
u0JvH/7ukJTqrxghkHUiHyjejnr2V9/Uismhhh5rKwMSaFNgABzIlpCu859+Y5FTUmES1nwzygxD
pF9Uws5GNDJMKScqvdnE0iklb8YtgOa8Di1Kh8BIj7/ucro9v7CGH51Ccf2RM6Xp0xi/3sy3VuZh
FezhU8ZoiSmkSVGTQ6+4+XllilOGSoOwVSyGf/bVSRnVAg0GOAjJ9d7kUOctJBa4rRuJC5bAtv1/
/a/rujVImb29oel+iFR8GjzOOzXaLbYnJbRC3RPR45sDGb9RFnBKIfX1WfyC46kDLRcX4pJh0ln8
dknJv1AvYtYeODZ+FjwgQ+wUXw5A7YB2o41BLEFRms3y0KSCJIuEzY5NZsBNMA5LXF6LLG6q1UGO
ZkUiMilNeDOyF/xu0mjcS75U1pybvBBvHYWJSop6Bd9G+AI8ObGKTKijK+cAP7Ei+gi3uqFOiKhl
pgc83d2l5Yk1rYxS4HpGVnHh8YfBYHXXkBTzlWw6cje6RzP8h526FS1XesuWM/qHCYtqbfbtCA+K
zul64LX/xyrkgkc1LE5IXGKSLI5MAvZcOZAQWGq7Dz2vC1lndjkSbNiDKp2TP2H5NXzGwqM2efXj
71kuHHO/iZHtRR4/c8DrfckJMwwho3hDkUhcFM9VsGWWigoqjyh6IYKKO4GrHrTZNLECFDon+6Mj
dJFxPSGtMs2dJmThsfuTlSqnBpWaiv3ZNp7po6ZLtwy2PQfdOnm9PCcifw9imqQOZiMA+w0RMciE
ZXTYrHlSXmr+InJURSGGYpd4f0T3WZHLGCgjjUt/v6mDbrioBZgznREMEm5iPlX/4ntSX2fanzEW
4YxIKzWNYbK0LmhICWwAL7QnSt8Y0uXOF0eTuS64Z1eVmi80amiMg9nGP42LXjsP4SCpmgH9ttMq
bAtEj+o+0a2N92Zlhd4H5Ioyhjlpg9IzXN+w7pKvyzqXis/bfS/DF/hz/verw9H4mMXw2aSpSxx7
9OS5QUi4mrA81farrPou3tHpwQCZdWZrrcUFZGOKEzGB6reijR1RJdT5nkp7fKchCd9/opDV+3wS
GkOA2rHO2k5ZxzKxe2O5ZKDKtcb/3yMXTorYvY1CvsIYVYBsg6uZnbubgOVjejHsU6F24n8y0rY4
APgSn2VMLSNBKmmp/16q7PNB5TWoBzCZKSwrjnkxPBWDcngRGMdnbjmPHXLSIT4U5UabkNjYKUlE
+VNCDgWL7zIMPZRvkWPxJz9b13RG7iZNl9SfJ/XIBzp2vcefxQoYzSwwkoHgWWjDmzP2x3HdTfCI
U2pynemR95LEVAFPjexyUUSTcFQhsgKwjlmg2IJlwQOWJeQgv9rgEhgKSw/XrRJ7VTMiIGTfUH4c
zh/wuBjHNkvmPmV/26ykseQUpA9UWSHaazaAFnUsB74BlMgmASqyEpfZcfD6FPnK4isSK4aEzbUe
8cw4dzjOXAU35DJJau219VukYN1rtkAtl/g+vh6k4z3mobttBT5A7CoHg1tYLkBgtVMV9XIueb5l
Wddfo2AGW93BWlZ4ELB+dGJt+iuv9ZVCm4x2SmnxRmgK/OOHqBJxnE9e5BQPRxb0RDxRDoiLjE/Z
v3C2VrIpOy5/E85j5//Tr6xOGgoa6dwL5DWbFfZYV9pBfEXXOIfFuzF/qXvi7BunbcgxcB3W8oy6
BcrgAz5fhNrUl317hgrn+9q7cSDh3mo3vLmWU4dpRgnq+EdY7R2ifwPhF19ysBrUxtzrNUZOVyms
hif0C6UXbUsuqD+7K7glgItbhDeLT7TH57pO/wdTpEYdxqlPnMGC0ewm8alX2H9NC9qO03i36wSh
e3ImpAcN8L2WGsV3Zx0zVI0PwhU4CYEcA1KzyBjte+FVajIvzgd7TO913DtgiQ3OdUdxy4I629je
nk9Q3sau/4AYoyLbo/s1+hdSX1AuuDJWC52RLD0zf3K40/UHOhCsjUuJrPyYx9y72iuWDv61k4AD
gYgEXpTMylpCj+l3LLlkKrX8GrygMj1ksjQBxXJJavR0XwgYzwxhHYrrAqkpP0pWB+uT6jvBd45e
knspDySzmL28GqNXbrere9o3Wy+LMP6DOPH/N8z1ytudXu18TnP/n03k+8QyuZs3lw3gYkA6rEqY
et6jyQB1ZwsCka3wYZMTkzJcs8vn2K2DfuUzhyNqAiQJGUyPFIKXvp7DEkALPUimVjHtlcFu5cBW
K4fRjJwa6b/xfb+UoGi5a1XT7SIurFkXhRGX5JKWB4lxEP/mvBEmSMQoqJJE1QkmiM5RaimDcxP1
r1jqd2W0geCGbbTgtG6YUOhMNTdULbVeLQFG1A46DvssVzaE79EzertSbT2b5mJe15xSjg7ps6yT
+GiKuQTPJHFPVweJzKgces7eVEaqGGYcQ9NvL5Jtfb0wz2yJZTD4FsKIDeFZB+PfwRl+rp5KMGuY
oWEwE15+w9rFS5PgZvoYF76+Wf2LvurPPwDyobiIQ9NRMY/qk8z4+geQz3rC/4wuFGgt2ZfaVJch
iXDpKOUl+QLQuzf16xcjRWAVDFMVjL1Wu1Dl9RtfvtHg57ue2P/WfIW3xKQwhjQVSARArHZjZHni
ZWMuFA7wIyVv6hQZrxu10K/4unKevdNM+LUklp9DJO0VVkpy5wDGd3PTd1Dw7nNnIGitr4R1APSF
JmkjZOzpn050W+udb5Pe9urP8to3op+vSm2gKK/99UYznROk6PDMO0ZA47QAkOrihf/Y6l9mTmOH
RJ90ZfHYxaqdLpYxSOziTDTc7dN4nxw+1kiRzevbNQtQmMi63Q9iBeitS88ypdaX2UJOX2S8SMSr
KvQhjfhnV/RM3I1k0poZWljQxfgciLSGLEpBAxG/TcMUEsqhdhaoU97RHCLH4U8dBjQX81Fm26Tu
yxZnWMfts8kEOojwj8g/Ui8q5UodNyFloLIlXYODAtTlHNA1DpbzarjeYFhxZRtnRPiiGJewbkhq
2tQddazua4AefZBb2mSjPuERg/9FFD5Syu6PY/DlnmvD0eGOY25gO0J5uZEF7XXrooCc/gQ2EUU7
8Fk6ZvfWFj+hir4GBlxcqmlhjKoMI/rxXUNQukR6Kx0QZm2ousD6pHxbaYdQBXEmDWUawLNETtQd
c0h/5N3+bV02f5XU1Cjka0iLt7dD0oQ2TrxVRg+yNBIL79/eZOa1sBeBbMW2dbdVeG8ETqNG5dVj
KCgUir5FW7KUPa4/Ye6sqW4GjOj1u/CXXnT71/S15gzWWVfK+XpQGHthOh9yYteCdyMQtSPNxc6N
jUyxpHc8Mk+s3GD4tCdYTlsMAGPrcpOUmlLYRav6p24pfBCvrNlljADnOXX3D10yOaXFwXrSAWeE
E0WJeJUej9lWuhkxCi4kxWQjfdP0W1n0b89ml9gJiaEeHwL8D4NfpC54FxSeTVxTm4qP/6cmla6y
J0tHUbB07JlqKzMd9dUlDwf+HaAEtzwz+xpiU+Y1A0BCHiLh60LhEyGGkPek+wceIuEBhX+AWBhv
w97Qdan+XcmkSgJtVRTlcyX24CWMO3/1iIB7FJob0209HdJQ44ECF6fPaEGzo6BN2fF32/ljmLwv
S/pnV/Zhmif6VnqRiy3Yi65qPO7SgXwjwycpdb9kO6fXiLNbxy9lMNXW/QY2qA2oC2/sB0sDNS7O
4TMitwngPDR9GIhK1vyrz4gF4fMiZRYxYu8e4RI5QlDY75hNSn9r5VvHvKcaVww4o+7aOO9wHjtt
6JYyUZNxGSPo/XYbtMRp5eID+3cMvEgXdloDqjp8tLJEdkhbZD6w4nvGfXKjSCKly1LS96oenoS+
aB852bJoezJD7uDcOP3tWGWL/M+bJdayT28hOo/mA/yLJei6rKrJJjffq34bKomycRGCIl9BtDk/
AKQx+Q0gXIClQZdAyE7hLSoKeJZolc/BW7PPUkm585FlzuSFAnYKOrkexbyhXcaT0cgjkIwmbhgS
Y0nPTBH/xQ9rLyGw5tqpSkxjfTBYW/r95IA5yZVDfPbZ839K6YP38gsJ2X7dXgibmnVWpuaYIPic
Ntm164JGnDPCC0GaaFnqnOQ7gN0aOA+SOeJ/mcHT/Ldzb8XxFcPOwRw/gOxcBYKIToJ+sBB4ItL0
JWtht33oZCOT2SAqxkSj0ruUZtrM7PxcTAy0/hLJfrNpuNeaDRuQUgLln2Tg7MVaFDU7e3nHsB2N
i3chzie6uhfHIbJmUL1gsdqfwNmkUMOpeRWSHQj68dUKuun4jzsuphdOdpsfmDwa48AeWTctpAZf
Z1sFJ/TRssRueJh9yc5BG1o3W8ohZCKvS9WTm04/wnRzimUjRPjGXG2BRGsnkBedXlbIvRhkbgbO
kYI5AfBdDxoGk+n3kvbMNostrwmypRAuyjjQ/Hf0J33685iyaKIQbXYXGbILqzPOUYR6gXUilBPD
1Fo5E0Rx1ptjRcUjcuome9fQ4OSc6Pvc18atAeAGmCYFCXR/mp1cZPdb2rj9Ey1zg+vIHh2P/rwd
6kZi1+HEV78W207/MGn/+X12fuyY8QhtIwNQc9vT79q/2vLLYIfEMdDooWJilS9Ndm00lbQyfxWG
PqQ1d2N/51A86yNti9QI2Lg0LhC9Kbft/polkplsxg0f/3R+fdOHLGb0sXMv/JAaEniDDfnZ55LS
hEU9qgouRE2+41Vaf1BZ6LOHVLJwRIiQJDoPg4pRPpHDkjJNxON74dXfJTxRMmQzeWJL9rHjwPKF
DZTqT3SoyNWnSnLwmXxY6SK74WCuM0Vkk4qM/nVC4VvuEO4tbcZvKLK0T7yM814sIr0Tw8HvhNIC
QFhruw1uasmoQnoOhKkk0Kv7Uoqd9NZqu+EwBkQOuGHDyMJnTQ8wpKSi/AnfZUjYjWdIrFGdHglH
mb+s2XHHpo91ZiOe3EdxCegg66HN6kVVoMgMp67+qTyH0s++H4sT0sa5k5lSUNW/PkOmHSxcURpQ
+bN7J1/9suZKOXAr4uOBYTfhwAPeFM+qnMQFZ5FP7Q56TaE4SyAT1Krnq09Af4t2/QCWTQuUAm9j
T4kBXOp6JZQNwWs5XZuBuRyX8n+wEruPLUKkxxfV/1ddKNf0PupK+cZpFDQaa3kPGLr/rXCWqCAg
ssiegPTF+1RcbJpf/hhXFGh6FmhtvWdtnW0zcQlE91HHUCfxIMq+yUrYpg/Zx51Xs0DXDa79NMfK
qz7SRG0QYxu1+39N/7MibJJGCyXVIZGXAFbEYcwB9TYaQvI/Zik7fe+VRIUiKsBtKWyaAY2lasgb
lNNCgtwiGNINyN4ZjOSf+wlm3r1NSbSsJXNTzd9OV92CAP9yCVp9MC3zYftLea8UyN9P/z/MtotI
XkzV+e1D2SyDbvBAurCW6T7UL3q65ps7K5i7bX48P9AFB9q52rcl7QdtifAMgZqISujtdKAOeIG0
czcUl9BoDrqJaESuah6dwqkfdwdIWy1piPEMmtqDe/dsUmcZpv5bfxnXMaetC+/v1pyw7uM7jX/g
/BPy0F/S+2gmyLVjyGg0MzWiHQutloVKqPgUpqctHMt/ZmV7cgwLFrmqHrlAYth18ERfYvUqMX4x
IIieBGH83cF9aYhS9AUZUt1RpIlU8kQRRH897OVvvjw87NYDbq6Q9eczGl02JraDhcigAlMYetHZ
u6nQPS+aN0xYc8DSqNHj1A8RQIDl9TPqYTUznUjJUF0O3InGsmAEe5BzHd36vLJTPD1qJdsq32l8
B+3tZpXuyU6n17d5WfQaUE+5lkn4rwXZOfCQw7WRoa1BM1XiDoe008TdqcRHDgvgsP/rhuV3NH3K
nvLja7uXaKDON2fnjSTZ4IOobv60yxwXMKMiFcvOuDlTyZBVPq07J7gyfTzGR/jyRtI+mfgUd091
YMbex0ZMMqn7SzvNELLZy4qiMVtaeQLNFtq0z1xWVH1Wz/GMY2EDHHvR3J9huoO6BJxSVKBT/UhJ
ZV/7BeAp5uCQIraXJdD+C2TzCkG7K6nZ7KY5okkFglLMT//LoCTnVFENH6CPmWroWP0YdF0NNYYp
dNdrXHxLZF2rnWvlzqmnsYEWwTWbJhCl7hh7OzFVIF+NH2d10Mhix9TmO8RHI00cP5dUkInsZ7ip
DJihbMa8KCALwXAemZ4Jh5vHoW/KpsDOKrt2AVdwHqA17BpQeSY+DGzzo9ydVpXCVFBlY6dWaodN
4dt2C1c+icpW8PT5qYKNuWJA1DoA697EpAWCOYGKF5OyeawF5lW0vSXdUSjggUVXNsTuPC5xsjJ3
y7AeFQhxn/QQQyrtwuRKVINPAPoyH0MrdqSbhtPPg2Xu0cn/XhVoCfNtNpbtA1z3WxdG1IwM70Jf
2D9w0+F4TRVtTB+w0fmIRAinSgChGk+U+vwTupu2ILJF2njpCT+fZd4DYtM567L+UPEL7bS30VgK
2DWB13GP920GxDo7VbRfHo+ZxcjmoC5hDwe4yUCbrFX1yLdyIAT75Q/+2okmPfGaT95T2CXn/Vuu
BRbHkBGd+ZpXJRVG7NY0sa4J7IjGLtEswvU5rq4rDavPcPgWQ8Fwa0VARHWlAik6l8jPENYuO18G
A8ee57I2BfRPN3GPeTkKQlZaf32J534XWfJgZnbs+DSD9O+ZnEcIOGUNdT79SWFaxtcJaVvRMvoS
KtA5nCZv6fSxuHC+sAztsRdcf+qwsD5FM9KfeK+xNjQ2B0cv4LdEeBSMSzrlz28eE0uG5xNH0l0L
lJFbAsklkOevIjw10rgeJNIUeKAwyfL2IVUNkV4Y2NCe2Vqt7BHo7tHE7wjYq2vkhiYxTbskHHVv
JJNxjWg8Pa78p+fZeoeXTwNF9QHbCN0t/Le+0XKet3Y/p6KiVXwU3aZofT3OjQzNM3DpokvjsLSn
ODTIlyGnKtepUeegSdaAd7GdChNj5vNHKJCkqf5HSPwipWilCmfZGfZ5rWiZjfDXzpJYqqIjv7Iw
iBS0Y4XOg99bLlu4T+Dks+fJP7Dzvp1h8yhtNoWXtkuxjDgVUQnk4z+hKx7edpLI0Wblg1Y904wU
/gmACM33vi9zbggujautCW1UbDG5FsAYNJNAo+QeXrX1pqs0zJ6rvAIwicZWfHk+n7rFduT33Hoa
bnGgEmS59oCgB7y3sz+MIrKMpr0fQ7rH3aDi4izwgP2RJ2NaHZuRsMWH+WafDlw/OFFBsTBGum+m
OnZEmQ/y29993fLwplVEyQGBJW9c+X00E36xDsOshuMeoEzj1+YlK8p5o7Cb9s7eeqw4IRNcBW0A
vKbUCd3LrIIDzmOQC+X6uXWRaSwPgX1xMrz74R1s1yKZ1ugOqcK2y6ZlQwXzzlEWMKS9D0CbKlok
vaSDS1nsoy7ptpsEzR9TWh0rQ+PC6GcZTl6cPGOC/5xLzT8pl6SV1I9GG8uiMNur3ato4Y0FYwYn
uAtTWWB3K/4bgHdk6NLht2so+WcUvma/udUBCJqukNjypfsCs45gr1wdT9erJHMiCQofK3J7iVYb
c12sWChtqegKvLj6L+CA6OsfFNUClk3ZavTRGcwQHqDOMaUMuG9q3Ooi2JgyY81HQVyAG3ylFbfE
uxXd67T8ov5F4yPrRvwBl+YU7J/9kqn0e08p6ijD//htW3RzISrNZX6SBmms8WxTT4SXkkw9qaQM
5wvLbaLAb7yDGA6uDb/++k2LmPHeYeLOcIS5iS8tGNn9EzZxQL09UTYKlbq1Rer1rn9wxiVP+9wA
eeXHMsqlh3tLvnf19BUZSHX5jDjVeTgu47i4sLO+b8/hy8EZCjnad7buq9ffxmy1gSoP9ni036Oq
tViGI2rjqLi0Xuz8hmxkRbJ9YrJl8HurigKupfQyiowFLHGa0B2UtARAq0H3mZr+htvTMv61yx9j
X63HOeUxixRGTzoWQhbSd876M0IjJCNYsh9R+/AGhSklWf5FqlPnM1u6V/TUEerUizpyi9LWPF1n
+DjtgoMyy4P6ZDY4RCtMKB3702r9cq5CIISbhUmOUNIvaF6lORYV5wIkUJJZNBCEN+fEMv5UWRnr
gJAsxZIDDWDz0fgO54m1bXp9mF6dC4huRKZcAYTuI4BoGEiqZrNumT8/944nkV9uqHYq4n7kdzKP
FYkHd3GMFLKLbNco7oEJoYJSt/U4mZYrdi/wDPbaLugYwEqGmLc8NggJ7nMprCzjHXwuXbz0cVtT
Va4hmlxuk+XTOthwLmVSid3wcWvaQ5sgD3DnVUTFZxaWLi3gJqdHXCJKCe31QQcO6XEA0k/QfjwR
0UvlNYIIhKmBhqXua3ADrHZ2MYjPUCZlg8BFsrzh2Ao+kResjyocEoIUwlufSWUVAC2MNLWqmvNz
DL2dwvBa2N4ynJrlgm6ennk8ElDzGHc4iFVp3E9cU+lUhqKJ/HHbdbZOJ/Pju6OMA7Jdhf2koH7A
ikPSv4JXq1XwLldbdhCw5kGBw8UXDLI9PqV9QUaQfEBnZpre+ViV7lNxOmy8nHADpNn94E7Ld9r9
93HmWx8vB02WWi4Wm9WNH4ajYCmWIxbnw7zXtnbqA0ej9Bc9sYC9CssmEJLQ559Rum0NOiNFNIQK
t/naelvK13CcHQbkT4nNG+qvZWS/g+t3IzNCzRV+9PkBP9aA0ZGGfnYumlXEtCCwPttSKjvjiQRm
7+sVh2QwmQH+stt7b4HkBIjvVafOvOVMV6HG+XMiWidufA/rn6/JmxBLrfXRRCn47NDmm/ZLBSkE
Zotc4sT1PfTW4ZO9K6t7Lv+SeqsxzPxZVlW6ImWzpsgWv09SBpd85j2J9VXHhvKIsRbY2OsfSJIM
hm2ez0ZpdxdQ2g8TIa6GKjeCOwO28MWLQ/3Ijb/EXLceyL7Tz4ltXLoccMJYO94aoa8RhA5P0m5k
m5p7fhw7wpNwFBPWsT907yGs395Q46CkZleLmgBZ1erwmprft2qfpw0upIPleUPtKEZifmuGSyy7
zClLpATiBljdecgEPgNv1lj95z4OFv0ff3frnu5pxTWLE2WuCTiLtz6vJXc5qxGUm3pF30r877oc
HmJEOaO8fJxHmH1uSQ1GT8utoW/gtfKtLzvjEgNNJq2FvbBVjqjvPz4JwhJCjb1ncxv9ndZNcOxS
nSkWzp0eSZRA2fAa3h34ON/Va8z7T2BE3kIuWsGUVSmRW2LXvSfssuDAX7DvVGlrBEFBe1FcRSKx
QolrIVyQYQyga7tkHwUWDNtYl8FxMEQgtBgBrsIlXZAUU8WfD8sWbNCjGQDmPPWpTkhoLqapAf9g
lxSYRN094z1hsqGHfu2mVJ0opZaupk78kdcQUGoUG/Jb6RjWDRdxGC5LIr7qPE7tYVDoKUlhH+pY
h9cQU+BZdAkuNP2iX31Q7f781yw+NtkBivMn4hw7c+kdtH2LpZ5YklNVH99IBfC/ZIX1Ro1pkBxp
iO8Q2yEMxq+goY9BMrPMuO3ugxYhDrXHh1jI9g6eDt42DwaKSa39XYikBbAcybgOxbXXuPFoTe5F
dn89L8chLXuZg3+qP19QPiU17zPkYLUJWb4kz2maDY3/5l3tliwonYHGeBFj5+mPQkMcARkWCebm
Z3+0v0/ZE+PF6aO5W8Lpdn399l7uvtlyoFLDfv11XmVMXB782qGexg8sJKvk+8JRAtV61VPlTjPU
rtr+DLb8dQjJjgzWq2Kh/HPTnD6rNmlSn4OoqgiOGXHcDntezH+o3mF8XCar+cvi6xzlr+nPecfR
DtZnThg1Qrcmd/I7isdf9NQHUSmFKe4gUgbXTsQ+GltZlFJ+HJyaQ8XoCg20opR37sJZCCTAnyro
gI+lTC07giCfk7dLRVhQaRfPrMZslpSRQsfvKLYx1vhU4kRDimaYCFQP8Nv14N584q4JJxzFrJDh
lBYwCYUusSGKpy03SqXfC5tI73t/NYaLkNJrFzTuUvKdms56goJn9gJPRtLHBrK9a3xlnXrZW0V3
uTLwxSKgBR/4Dg+e+MAJL4dkgg0zgY6/5kdep6eo//Lf5WwCBNT6ojGs/CELj8Zswxu6CoGKOf5a
GL0BrW2f4wFwqrqAl0BwlpgzlnsIGarK3uDezXOprlCAf1BixfZrLiRoAqWc4RZx3RfU1hyuN6V8
C14gegkdQNhtzuAnUQDUwWhqXj0sZZroGbQO/bmC0cAjzjZ6impX8t6YH2g3nAwd7lVrF3VsJ3w6
79MuKYw7ba/lj2eLFHKrOKlfUmIBnRKwyERpMBYJukWQzvfhGiNY/zxhy2HIFV+s6XRzh3NQ4JbH
n35qaY7eVZgwrQVLa/oEAZVbobP+79To8wblOqQkofOPjJ2ZjLYCPdmqL46uExP4S0QtwuABzL9S
DSZy8nr1L3Gy/7gbyns+ZhGh4Zvlo9h/z8PofS1EHZ1EBMvalnJ+6Jt72OMkGjsAiTEUOW7HUJy4
LEgMr1bq0P/U8OmWLFtQSG4roGqX7ZuO9yriFWV9VR7BWCxWC/6mxyve9BGSkltwDPlNlmjFPQ/m
9mRdY6vyuSktzLWUhXhA2E1vY9QUHWMoApkabNbtUz4XeAW5bVp9aWkrOgq079Vm10+aE2j2s5pN
+8EMvjJbG+m6OciGHL25FcTiDfFtlfVbH/5Ekj1IH4tqetc2r7yiopynREv4TprMulMfxjapVUrk
NyLgBKXQEwqWENWFBZ0ddZgnwWt0Dxci3vgQUJ5wBcwXrML658ku8Yjb8n4gSOxVqXNBRItxqpq5
itapzNnENPHf8UUUBzy155qdOn6LEffvBFs6bmNYeUcUvql4USumjgjDfUIgo/wY3gdAaURt46Kn
yGyClQ9iB7KmfJh3GZjUW60l7X42iF/+VuG+7vFK6Rbf6vJLVZphpEVxbbxYpYHR61ZPSfSt4/E0
DUG8jzwNp28Do81tLTjwuQ997d4CgbUZ4osnIpRMvJd0nND8uri0sMDRUJ/Oh6roUHNYFeB27v+5
8ihtAESmhz5znmDiDyXBE4at6INynnbDMrrfw8IKu4XyuKLkOeja2/nL6CtOjLK3EUtui0b7PtVr
3ok7JKMSr59sCaOdXrWfNsXGC5VXXdrpDT9OdUcqRmgDdDuo/x6nmRPAswD2OnXw0OWGlKY6ExTU
EyCaQGz8lmgQ3jCIdg7OQ4brUacgFQg4rvk3GYYRN5q+IeMsvbD1367hYIdpuoQryZd7yp7woP3d
1Vv1EdoSTIWgP+AaVUgIBPPjrcL5UhpDbZcv9jrcQ11D4aCNDOByPHz0A8asDi/A4u4bUc9LlQDg
V5C0eGx/xq7eJB6blMQbVHWoQr3zfOrym8zNtGpEJv8vU1uoFFPF88U5sKIuwNQ3dwAdB+Lg0m8U
NyCPCUk8olPoDZI2LaxhtCU6t16xcU4s0Muc4F0x7ygK44UBt1VFddl7RRsvHyOQZDnFj/SEWYks
PaO6BczpBuBq5ciB+tJclBOqrDNLUep8a9hwoPLoTCwdyjjcJDRjqZMw0a9UIDEdvaKKev9JQEXE
t8eL9gYqC8WT4BzdhxpbDk1rv0a96BZvE0joNUL0mjEvX89jt6D1daVxxhcKjzFDWI3qFuXAb2dG
Z/XFddRXwUYxAWBtNmrjLWLH4IADb5zaYUZl6v8V8964/BZG/GMA+r9Kc34UWrbr1xjBiS3wK/E1
TnRJHHmjXOIXNl4uMkHCgsz/sZTBrqLkkzJ3uiaW+ynM18Qb9GsVGoqO5kbbB3KGqgUNFhz6vzMm
JtnBtZcWpoljdiTqAd6P9+yXu1Y+xwNC5NsN97jlb5SyqR9sAQ9Y2Kk5LxJond9JsZpQt5aza6wL
1pGzOl+g4rljj+ZPZJWrIpCKIgm/8BzeuC2VdtSYRYClJnZZ0myr1KZrKjYqnIDoZvDBpEbSzVK6
kwrrxF2Z+VK5/tNshad42c1lsejoQvHq6DFLV2LCOZyOSo1/mx+QVn4pivmFEQNIBGT0MUyacg6P
GIgnddCvq/jnAtc1Bw4DK9ugwlQOv0CoV4HJZs/T2cI+3f8ouAJx67+zPRZtAuay/36FFxkFY5N0
NY6egBDcLDMD2JyAA/uAxGnY7Z06LsDAax/voWSsXjZVSlMfhRbORwhFJ2C9jgtfpFcLclEnb+AH
rh0spspatQ3CJuU533SUSKwzFNc1U3l5KriO8VbRIYk2ussOgvSxnrIaKMdbsyV+Lz4uTu30UkN8
eJSCy93a0sFeu86lyJDb8oEjZhMcYL0eub2xV8E2tVPrKryl/YqdevNTJUoUg+BacFbRjqr5UOg7
k2QcFYd2thmMMYT2tXUKzFHdd9ogm7dAL+gGB2QWLHCIkHhatzT4878KibSB3IsWkjD58LhrqBGh
sUUyhW6/DzjJW5DtEsywmEg9gsPfQxNIWwgp8YbOREMrC2lpIqXgOYiZJkLBM2ZWqMWJ08lJF7qc
21aYygFYrniSoCv4BIQRmv1WY9hIcdowiNVXEYss0q/a4CeqLYSuoaGRqbmO5vbC2JUempYRHz6e
cn5BprJtmzrtd4RQTgh8e9ZIfet9LFfxSvK/dnSXDN2AwgihnRKv+yV+5H0MCq8OSbnpoDUSuSBr
R9frnYNOsA21qvjkE1Ci3HbdlXREtTWBACqxGb+1YHl6p7RCzDP4jengP3xhlrQ1yKKd9rZWeFIZ
bGY8jNWyZKImIj1r9+GzeqmEhDv937354iPnwi42fd1mb9i+Uzw8uUFw+oYBbDK4HFzg/iX9sMA0
L7vEb6H81XK4qKNjJ3dShFqqw4yjFR8I5vw4tv9Q3g3o+kgQUKSnFT5nmTxeXC53ifwrcCIJjCXy
CfWM0RgT9RparYSCCM3KZdGyBYcFKC6qIjgEVC5Hv/ySYaVzjhaebUC4B6c+wuWum6MQL7YmLrrf
I43+gistNWQKuSW6dMetQs7opIsG++rnAydkPwyH+NQ1Xt6jNMLTRb/gr9EFnvpbhFGmD7lLzLCS
V5nCzWn7bu224TkCqQ2/YMagGdBRwWkmLWzqBiDh4c70vsp6YPO+02lazGbaQaqclCoAURFMevnc
NFdhS/cKjCh8BT44arXGFZbCjlDn5z9txDPscfHmTmHTOeWU5A7cTnpUmZpYqqTrxWnuGbHb2u4f
Xamjk+Qm92V95FVKRcAFqobY1aHNysuMJox44MIOhmJ07m5rqqCUJ6VxVoBTDSGFe6m8CAgXlsIK
6h3FVXqkJNneJKJesB89dHCal3X9cyXnCQ8aZeXkscJE5I/iLtw/dkduhg1g89DUIG4MeWwsfwSD
FUKLdzpBW1XW1DWdC3SDiCHwUl5pwfuLcbsD5yiMtFMLRxJ9aJEQjd4SSXFwN/Fqzv2ujeHYDbZW
/xKzQjZied6R9tBuQ9Xw35BiZE0H2/Nbwp1ROn/cLTnRQ39hz7SY1JDvB5tp+a0Xrdf2EHct7tFj
hrEI2hp7BeVWCAsyGb5lbTLS1oKFgfP+Xs5bk68odvHykD9hlfqHUfkCR6Zal98CO8I1LMMqM7Np
5Vqrri3kxwrDrWoyVAuwivbow/+6ZV6G9etLLbe7BxSSSDHGCV7csobdd6eWrLVj65SVG5LpUbjF
MuErp+1uyZNUU/bt47ymJFvMrK8KdQF0TJ76Ma9dlimb1OUdonh270fYAYIlctlQ83cz0BVwC51j
cco8QS8hwRs5uqdad1CilntMZswVizC0Ykzpp/OGHxsFWJpZNnFJomUjTwRnauyHK5stCDyskhdL
2WdBUsRT4n2EpQcdSC181ix/PAZiXfLK8LL9G+LxWG12pdH1DnSQM3t8Vf7cWDnOQ+XoJSfapt0N
cmqZ7ZCHiYJnTVoWtpnShSSSZJ3H+2mpje0C8E2DAjslx1sh1xz1dj1haLAMKCHDmQE5Ek9/RqHP
CyGIM/Tc+w+bo1sorBpcj+uPJ9AoSoDy5+6FczmPAfMzvGEybnGW2WEKpND8sEcHdNEmhBE6/Ep8
3p9SbSICkmtGedUUizq3Hval0N4hdgcVDltw/rC9yTp/1Mf3909xCfk9Wb6ovT/nMvfIgj8A1PLE
PreedV0UYZaa3Y7NssACF/MCmPvVNsarlNKu5UErH2YK7vCjaSBpG7Bpvsn+oqdS0QNiWA4k/V0m
CRWKTUU9vAr7JVfa54lqWPCol3cJmllWBU7yHWVNdryLl8a0TKWLyE6cLPpNZ3JaDdN9sPgbYop5
fRlOAau+RUDElwPUhKIzSu4/Ean0FBnyj9AnDogILnUcU72VJjbpCRtHOGsWYhmAQ6ojJ1h9EQjy
d8TKRrHcMzdsa1z0RaGYnmjR+8fvIIwiyp9mDo/o5FyzQdG5W9ldJE5XvY3sR0tlvdo3GxGvMP+e
ghO7Zyk2tNLqT39vsamf/7tLIvC+kglDJurZCFfzOqaTKfebP+O7a+OO9UfhWDk1B0xbehxADeny
21LLpVRnZqwM3XY5U1aW8slxje0VUDM46K5X7xAcfzAOtcLzrpF8bZb15/i8OD9/vEcOo40TOaS0
XG8UyV05K2RU9iDkvES2FHrOpbqLs0XTi7UD6woWH76xvm/54YW/w3Bf8URuo7Zpu1YL3sZaQtuR
ZDyETbSNfUKffqPL+oeM846OpWB2oU+Hbb5easX+lSrrwhrZLxeROJTR6UgxN2XotYKzUkhIZ8kV
9JwhzYJ0d/fInO+T9oXdUZCpZOGh+fD+E1W9fipEt8CkDHotRe5XiIvKApxJo5yRRtd+9xbFAlAc
eM9/G5L6TAv7zdkN16sOR4QXZgK7ui0NvvqPhiKb5wnibqkCP3phGt4ECnMp52Xf/Mm6LtDl/bvI
CKaMKEL5m/IEXt9hk+rWZLlwY+0ybAB32lBb++VaM9S0QdZa09PnukVOKcOUAxKLZ9EP870hgmDv
zAiox4tHg9h57dk+r5BErWhajJQTUNFDuLy3iIsF3IXz/+xmSDVHhybMYA5UgGHXJtxFfT2NSWdC
0sq5oXHhg8KQqkLx37Yj/yC7+URtoMB3uEB9Qkya+M3lRLPTmQvosd4LEBQi3m0zRmPKWxOSsfJR
B/In1JAC9jDmmRPLlnY2FO7fdtSu/pq6hPvcqjS2lbrLqXwAInpwRdnkthEakifsKwmZvhdYdbge
qzPOklZuTXrpb4DJrNfEjhlsABLt/Dl3D2oV/s8pdmTe8f+QrwlCcX5tW8nUjy+OpZs4fD1INXaS
M1+IXEoOhwTYTbalLQAg3hlAw0ThdJxCs+UAHI/9oO8Yr5RwUGpu9/XYoPGA+UeyVYS1EemQKD55
ZrDlEkHs+fCT7F2pRKbW2PW6GYtRs8EL+dS5Dj0bObxZIzpZCzSEr7j+GHq3P/hUtXQsnnENXNAN
n3unW1ZNHB6fhStfXBToKBy9eVA1RN45vWQOLmIINpr5kgmSvnDYY/G1f/sojmt5Uft9kV5Bvqii
AFJ2sLm962laYf7NhKXU+2fTqtB5/F1kJbZDjaSyKBB7QUVdLBYnzKVIO0wn7zEQQVSpu8Yf8Zx5
A+PtnifIDlF6SJMnAPuroXPxrOVmOdcrpa0M3x5DMC84QosTRIeabyvxzhhUNmKceDbW1wP55CH4
3bUXVIdBD09CL/yV9LSC+VUwxZmCLF/R9iha3eDAQxG7MPRVIWrz/9AAoqrOC9ua193KqB1qcfai
mr1AXL/p8o+ep4Xw8T5g8ec3Bj7MXxOtZzhohKitWE6oF4dVN31SHdPHxO9GWi3FPtfkfEZ43DCG
MVmbW/DD8nmDgTkbdWhPg9c5OIDmDCWquGYe5LMWV5737VNhDY/WNJfVRSCLMiH24SefyyM5XWrj
oA0s4ijZxsxUCEAFxt09Dgc5QShkanTfnesBPoFJra5+hapSzxvKHuFw9jHUHJtbw3MUNUr/YX7g
fT6VSt6GnFgawva8OltCVGKG7essgjsN5tjaMnr2xZdxsC24mnx0c7Wrigh3/SGFjX0irkW73nL+
Vnzq1qS90Xog7NSFplsMISk71WECm+SQNwfpEatybjIB/4Vf7aqhwJ+yTZVhMgUhh1LGNwt+6qWg
HYb3uA7AwnhLB6R8VkCqDAJDvpeXHXAkP6P3417Dsi5uQw/BjgjqreImv4Wcb47Fsv9f7qplwmep
c5X7mJTggkR3NZflM/ubqFilChIXYXGv5MbSroRzY+F6r7qMrV9xjTgs/pA1hPesOk1a01IZWUCO
1vBNxDJVr/+4zymq8fz31sGtAFry6qlg1gef54g3vaiaE/q8Bgmk2lLtfIsL1MWx5bKP6He01eKP
rKRPY8b1A226dFlQlK6vOIFQLk6g/gmJWWFfYh0HhWjRp7fHTLZYxAh0t1YWGq3RKPYFzwsiip6i
J7kQCASv6RVwFAkmHPHVhMHIT2LXO8f8JBoaqSdU4xK8maRV4LdXiRqRYGkGqZDCKXHd58lIHaGP
xOYgRcFxKnKRiY0Coe8Qs914ieFq7TCwz5tb7X58Qv4fEN++naOSnxxQ5gi4MaML4NYtlRvTAPOA
TJnFb2pBG2NE9/aoQKTTojcOqIC6aJwH+g223rf/bhosnhLJyT9x3CliWGn499XAGC+ZBK5ZIy0W
O7HdpHrovO5Z58dOFnGcTOhpDjXSI9p2o0+ASY/I6lF0ofenPC+DFfyPv7dgZsYW80L39rHAXrKP
Cr+ycZIZDM1yQlUW0PZcf9IDFe3Qi9chkLlvNBM5hggc2tlD5+5VS7/3dGTHz7kVinFhLDfxAg3a
O9aTtZTxK1UUy9fQ9wLWSIbbZt4Xd67RfmX1OV7mJbR3MFYeBDdYH5nCyV80OUSeBpQIozm4jHq7
a1kpQc2CFTkg7dNHNBbQJy6o29bac7QnpT1v4l4Ynsbu72mLcL5HmLh1zEVlzRMIaCUrittYmUjy
lsIOjHTf5JG93Wlgxf75J2mGFlRMF4WQk5NzJFDMg0Aw+olT6PpCyYrz58WU/3tXWcPgJv42wNtv
Jyrvd7+J7aU91ux47z6VG0TT4c56c1U16990lpnHXRo9J4cTTGrNB5/j7L1L7CenE0GPennAFrFR
YraUNO1LOLYp0g9+DFowQB1y9FJmKV+9B0pOXsf9M+NiY+hhuBbFf/XWJTUPdz03dh5oOqF6nmdV
fV5eOnjwvnU0h1tUlrrm8J9h6IGDlWMSMw0YAbXla1xMrt5By1DPKqp1uFh1XIlLHOL4kBYNIC27
DVRyzNLUGo1zQaDeYF45DkzjfHlS8zoaexLka13b9X2SL4QyMf7q7KR9LUHOHfhA0gv3zX10UN+O
ZB/MNHgWOXKrrMz/BmOxr4N5SekK9deERNge5rgz5TcyvpTrwFPI0SM7Fs7pE0jAIp6CZtH78PvA
Ni4w3KseDkjzHW6y/eFPU0zK7ZzCOgFhSQelIE0v13DjkwPfPwo7QscanZFnCeFuZ569o/9Oo+hP
QCoWCaBGcNlxjKTGICNhdcdkIhuPRoaZEYAV5tibps3h5Z+MUvk5I4Hp1K5KRTqx54FW84hwIerg
3wTJ5ojdpoC/RmEEt+NQ256p6mxAwIpDwOXDRVGMbufhZU9p4cjKJM32toSHc2lMdyVVpm4KWXio
U7N6pT104QvvY7YlKAKlPzd2zU1QcXbqnKaHTN+Vv0cd+twmeFQ+zzF/RbEuaDgCDMd3RRnwFYED
NnakvbtJtfOShiiMlxjJ8YFXEKR1QZc2tLUMoGV9V47FAlFT63gqiMxIhuE7jmdGy9bV84mYoGng
NgIXuvw1TyilwZG/B2NKAts+9O/8DSsSN4zuAORX4FALnKnD9wiusotto86nzf6FQ+bybuCAol3p
S7RvHkBp4S1elNM40klnE4hIRs98bqznxVns2vaT7AjXbYrgwUHwsP3FpXDKCbD4L+8CmYSJxCiP
Prac1/lCC7Z6rzZgvqku1Wcg4h53vxYDkyEXp9FA1YbMfDCVt++EhgRBQhR2i9Ew9PEs0Rd+yMT/
dq0NYwk5XO4NQBVR6Z55c3ppc6rxKi+aOo/q0OzDGcyQXundMp3bOeoFFcQmuET3/WaW++2ag5gu
R4TpnRrQNP5zUyD2ADXPvCL95vuS9yl7vyOxU5+keT1ucVRb02yVo2cuciFIGV2g8O5BN+ckXO9z
UiNjN/I+aXs4Vum8No8/dTx3MV/JRdzQQoh0dRmj3p/kwnZlUtjoc1DzEBMXoYJw/0d+pGmWFV30
PfCY+igWQYfdL1D9xdup7NeV9KS/NbXUEFV+wE3QmbXsbuwx062Lig8cj1VZNKG9KSDM22YcA3YZ
Kek5MsHeDQrlNZVYiDQ8JSo5+/4GyBbC+8ySRIkOSfQHYQwKJbQDys9VZ4pVB6Nar4k1U4X7s+rl
jP0pIuNdnwPrzYt6426hooUVs51Z/+inQjOJJ0kpyGzjopLg+5yN7PiXCNOTntDrKHu5eAckPXOO
zBlX+PV0LZ600RxfRSaeHev9nU2uXPxp9YnUZi1Y4NLy0qw+QAlT+ZCwzMtnOONqtFA5BkNOnUbM
4VMAlEh8uwMi9D1qoJCub2gviEu0rs0gzIK1gYJTDQrTrP0BuvON9lhjsfswSjtId6w5FsPM6spZ
/Q7Ybl8iMVAhxV37N2hOLfcHDcRLiaD9tYIkLlqvsKXLvS95w/80nPfF0Rvc+CB1FaHSAbYKRSBr
TYChqyc/xpY9nsJdSqVVuDo/+qTcdquNNFyKmzFY76tHSnSdEaClXwRNDugdQATlIs0kUfFty2I0
ruO5djxxL5LDVgjCfa1mF0kQ+DqbakFvR6bE4s6zdWJbab2Lp/S7lbyrIV0bwoJWgiq24edTtzB1
t2q9ukMqB2Pvn/d2XQn+kESiAO+byT5bYFYKHnaCe+8DeOJ+fTgufU/zswDSfj58cI3BOti90M+5
OKdOmmk6XvpFIegpEJm3aROZsYcbDUxaB/yUOuUE+Mdlnz8vgSiwVmxvZE7TMNIh059NECakBY41
JKYjtU6dsLiJrS/7pcP7KP+aU7lntukjTmErhAJga/NhwMXwH2WZOU+19bF3E809sfw+G3HPLXPg
ujwjTfR4hzJQcyaAmV2BEsE9yop7i7QqqT8mLdSFSIVSpU7+EZs4WcK/qHvy6pRbPkDEh4Nmv2ZU
/ZJUyOooWBffVKTmfBiFLO+RV1w3J1jmq2muk2B8EVVwqXZvTc1trCzn2q0tS09W5YWb/9cfM38e
D1px6F1oE/pX7IuZ48xBfSjnvtZlnMdGygSlt75SspbmHRzInQwxJzzGABY1PwuhUkZ1iKYDM++i
Igyzx79lP5vxP7uPd9r68NkY91qKZqoFOoo43LUyxp5+HPDdy+qcjPdoMhY+lKS7AICcya0Lgnf2
IyCp7Kr4Wd73OVOu2nraIDdOKN8bnbe3u3ulGN+kyewLKHH6/8SCTiReJbPiPrU4FWmQnR47kDLN
fThtZHMJfSOG+yz5Wa6H3JEIBzQUpfKbMjKt8xOwaakW0z3Dc+sOp9NFJxMdBzU6QIf3Np4qpOFc
N44NKS9F9lCGPErRcu+tR/z4jJ/ZseonwxZjMrvGQe0IWiTEM9vBvKE2pgbf8VeoJOAzR/2F8Py6
5zPcbDO+HhehKkeZkqGoI/TEcwuUIjFul5cymJqUPPrOp5+PMcbcnqNzdfvbLRf3xpeKdJ6JQHnq
bZUI5BTgF9B55Bv2D2TamEyXgtcH8+ekJjieJ04Waj6Pr2kYOFFr74i2D3B1MXDALzt1d28IkfMk
LZNyHhGYBx/RrSB6y6dcaiDIjFd6e0m+D+wcVO7a3NFGS/S9LJV3rPidOpNYNFTePZUmkYzbcCOj
gVjgU+COOvqIxzaOMRgHcOVt9J9sA6qhiFznpgKTOeRjfqBiT1OkAhy0DQTDZlJr6Y/8SvWAJttz
BVZxRfRCuKwKlQPKA7p/Wsfm8NVhR8D6q782q89ZWCt3oksRCxsryMkRs2WofHT7PZjr6Ka/8umD
GpwH68Y6O+l+mNEgFDFXZBMG3C7FPUb0F0oRVvx7eETtbIy4p8xaL/zdevQmAaTdSd/go1YJEDvp
3il5ff966OFk51PlMZq7SV/JdKggGpUtXsV26Z2S/p8RzBloI88g2I7w9DS03VuLlah6e0BQUTpr
apL5CW6Qpy3hFXodl1WGMhqSFFc6G18diwMNU7Vmo4oxLnaNHpmAs687yOIxZmvfhkW3bc35Xdm9
M1agFAd4Gophu4xjDNJUzs+vJlwLO0rpLVJWnOaps5S0qtSFVpC7fP+Ohp1FADXrSVqZvpq8itHC
IIy6EkOOUyxnuhA1W2aEsTGfQuyyf80ivSIDux8bOfoYl1l3dhstH5gGkigXLWULHyUcb2+CfCHL
xEjcrbSsk2qwvo6bdYIVPCT9e84S7yIGEnZEf2Rmw/kmsPSLsqOEw931rWFke051rSAAgJcC1/Ce
e+5POYGjtbcELB8/D9h3aVw+X6ZT41tIJkOfXUlT/rhG4gEjhKb7BDAP2ObrzS5pnWJtQ82kIZ8P
nfhja+WDAfuXSipwgmayRKfdjGor3JqVpQ0P0PQtcqo9BM2pTi9YbEuM/Z5HJAYlCFigL50qVd5X
PvwCRvLHb1I0uHzz9qWcuF4clCbcvB40IFd2ePIEgTXEdAKbAYY26/+JePXt2kedj//stfog9Byc
V7MPCNRjehtRWyUMwXDzhQyfVN9UnYPCJFTS0bWz0uJBuURr4/fY3ceH7lMwSQ3N8yUYyQX2eYSM
038p3ejTh6x2WwXJdoStrymrrrAxtumVtT1/U5d1cA/MKEEnpXWZ6HlFU87xiq8+bV+mSMdC2cpT
0SQjBJdFwAEuexhXpF/sEfa1DRsayg77Yt0OjZZvrUc0LJACiQdyjKPVVOjE/wyNKDdrguImz1fL
yGQO0evXfX39bfGHtx+ymVRUS6HmkxpBAnqFNOVyjrhinqBDpuNBPYG3Zi/Y434/1KoXaYChLwXb
MYgTlTunyyQrvA3tXhIHSFZ0yYdrqatal/UEwY5rNk8ph/dJnAtWEISiq3tuh7QvDK7rXg5MSgbx
h3PAlPW3CUoB7fRNFALBcEPxuH5xmL2bZDfug2TeUAEwAs18U/6OxtQEBN4k3SX5NeCzh/c9C2IT
4rJr0Urr9eb35EypIUmezq8/ikwldLhGW0cNBi6Efp06D4lI/T/6OcBnrXo14fi2atUiUnQeo8Fd
rxXrNlfKcQVAaQQgZpZy7KTmON19Fcen2sxSWIiLf40vrGK5cmhPNTuVCxqZ4bupGfwvBs08K0uG
NkYC26jL2/rs9f79WBGnsCuqyQQreWm7szsCkfvmLrPaP71k4IW/CXzD6RYqQxqjvrnLSHTkPHRN
biHLfFJuLZB1OEInav+UyZ7BWUBmTrBSE8TotmR1LLQ36fuh+MB8CweWe7btHmahGk7y32E4rvDL
jMmM0o7tInn2svqVbI5GeP2mILjhWVQ1vqdg8WT8lRATfL4KLcMF+WA0szOYv7Hi1GREYuufhyi6
f8N1KWiPJPMxzbuAMOTw2T1mSbqE4lmiOvWkZPoO8+ITqhJYpOV96Ie+JaMMIsRRJeBa+xBnkwsP
N4MC+K43Yldr3oDgQYfJ6r6Z/WrB8+Qes5PLQt8cWWtprS8F7c7UT8xeflX4LQJtrVP0nPgSCw2D
QMosxWTy2lT/4RGuSI9TX6Qxn7vQatqj9VwTe6Gvg0Dab+kSE8iw6VKajwR1KzhNEKXTvc7buTr+
WhQIPQHzNLl9Hdo3PkJj5RI5/k3RPzictWTgu0n8ExoJRAKHYGSb3WewPtU7IjuZXySzYyrRsfRD
Bp3fUYmAZLPfnvtLZY5nf6m/hGbTZTP3WrS1phy5qe1pzs7diYXszooekpdc6bPFyIIXAoafd7E8
QXB/XLrWEoy+MlyfGRb7bPvQDIZJjgDOgJwGkeCT+HXagbvRATN1eVwBeLG5nC8HsvNh9cZgC+Yp
6IdYlSCQucc6j3oUjrGSzho4drOVdFJj4KW9FXR+tkYbORom6h+2ClJg5Z5dckysJ+dcCAG54+VB
BnB8RUled1IJgkuLIuYeNSA0qEApLgP/X6bGgWM6I+dhVjvyn4N9HbYCtXafA/mp7sXYJhK4DHXJ
mzqT9599y9s7eWIlbFZA/+IY+nGE5CE7I2a/Q1upZKzCFgRgX7vqq8g6UG90ZGhHwkaSsOB1+FiA
l417MLLgKEWg9mLeacPpfElljXz28n10eWFmNT8kDlWdJvOX0l0VMTxej14ff5AvjQUAqJUeZz7Y
X1MyYxibVzhULTCojEuwKE+ltG+sxxmBvWITwXVCtIXAGz/y9x22hnCL+dTX0Aalq2VCqTJDoskB
tO7I3Yhe8Wcijxs2Y3gCf1BJzrjPsDPe5nbJhB0FQ5hoRPc4VnHclDlGQiWX8ZIL7lUmW+lPF2aH
GVPAq4B4swXxWplhsdiWsaGxqSSCn25hbjg+xXs/QgiHnTWl4Zyl4QA21pGeZRYIoEqDI6EWorLA
f+Fc5td/xWtYzkj6g9Ryj8sotibtagE8B1Tiw7g=
`protect end_protected
