-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
B03G8bYUnGQgjcm0xTEqjzf2ZA/vyOJoPcD+YQlt8ItYQkSVHQMSm6isfE31EH/cmZ71H8nZhvjV
+yyTKBy7AVKm+YMciGwoosbiOHx1UZYtb2vj0kIi5CU3kCLmvL451RKJM0oMeR5P1WTrS5YM61f9
jYAkoDsxh+g7xBLL7NZ4VarSrLKsHki7HPAcaaiJCh7ETPQm5kI2skPB5zycMJCnQUyXtePX1l3d
JOEsB+TaUmSm8CL1wQ0Bj67gknoPQtHXQ/a0IJs6yS0UiOmHYSmlPouZfIqDtK/fN/Hkun68cZMi
u6JSZmeIoCxXr2loVKgSPrzOwrMkzOFQozic6A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 24704)
`protect data_block
Yuj43Fe+ifGL3UQZ1Cyr7BIv1/uWMuR4WhyAoq0UWDeEeHsinhls3ahwPRF5V/Nzpi5eQZlVdIxV
FIxumDCNTFNAVxVi1Gt09zF5mUs6xPwb+Oj8BiwdkJLE88ZGwNw31n2faYMz7a9faG+HE2ggxu/B
ZjEbJ68BYPzM1sHq/9+xm6ky3r32M/moL3+28/8EDuxdp/MExxdK0oZawlHgjwupL988Ba5UglBu
b1tJ222vpIE5dlJLXyRbCTlvBeY7/uMUk7YJ4o8yyLUn9nyGS3iTtFF3KxtUxrn/A5YDqa8SXq8o
2U2/3RbhI/KbTeZuNZujGQ8TPKn1y4wJzAV1sVKnLBHkDz9nXfQO7vniTlVN1//lx3j1JdkYYr4j
1i29XZBTkHpyBeMy1rB6KhKeqboGhDo+gcTtPKg5lrD9J7pWcFzcQ/Ov2CYYNX+MNqJt7aFrAYoT
PyysrI66io+a1YeUSbpjkpLCHVXDta1ZXFL8FUsIFpapFb//J5l9up0702Cx9C5jByGWZc9Ufz9E
9ERY5uWJdEM65y92PC5bCITOvhZpcqes+5CLZxfW4y/3i5hzxq1shwobdktX1FQ8mRs51kbzCxGQ
mTAc5NU/oWo28cySfFmGoNhxM9rSmwBGsNNo65z9yOBzgtcNp1qnMNd4skZK6/1ZxYqorkvOd/Mg
iYm8dwpzTgixJ9xQajn3VC4rfWiMKbiJeBXxTK2STuXk6j+qUvCK4X33wUpxhZMcoN0Q6Tq/0HEI
EpsKqtzSzhKr6cBSE3x3i7Xseh0CavBtBG7llWjAJ03AJ+wPvOK3ySzOQ2wl97syxisVqlk7M1Rr
363+UEAPubYrSmPKHEvTL8787AlvqZdAW9wvXLq1Wl79K8McNBqwLVE2m0jzLtiGI1ILqTW3v9+m
Xvnd7F7ZXboZ4//HhP5xLiCMUl50ihl0PeoTFpaS0lGctMWxfCNJ2DeGcmHg4kcEgBF9TAvbiEQd
WodqjZ8gXXon0Z8VCCTDSv8ILFii5MVkzxcm67sdsCYwsktSofdfc7R37+TRrSl7QWOgSGehh+zJ
FRnhtLILb3kMt32RuOKN8SbjULy8Kjv7UOy8DF3/kyc0JMwYfJGhZ0/PQ0wBy7FUJd2xTrKZF4xC
VKtajXyuzH6S93JcphBhyFkBJNHbQ0fb4StKSGKvYLd84WUOpbQnJzJn6dtdZ2J4qYIePHAkDONy
IpTsDn1xQz/C/h/Si8jLfQrTiDHi60NLamdNq9Wk1h66kO9OedEREXIoLRG6E51xIxncYzlTVkvr
HJIhUpYdqF2KTzoPDWah5OSBONgdOU2TQHjkKVaJflxKQzJXVDrqV0GvHRO4kQzgp3dnyUFWPVEf
mGNlobWYYEV+G+NsUKTJyQvmcLueR+CzB6Xf3kCel94XabgVF5Zeg/qwptu/M+DJRNS44ld86C/A
lyUN0GSyKdg3AQMRZNVcgoM7Ne1RiGzpsgBhqdJQH7IE5uTBloTk9qREhQiYILn/51zp4NDx/vAG
I07nV1bSRbCeLbdBqkg6xz+5ZnowEToyUJy9JQ7q2q250sgkTOBJmO/CWZGxUHh58bA8YYJscDIM
bmK3tSy63zmG2hdnlN25HFmrqhObEPj1ftdj7pwXmQBGpNEYfQ5ElGGuJlYBRmXRr0brgDW+r2vX
W0QlEGBj2jbvdwtTPK4khkEvGRj1TCzTuNAitIScwHPyuWD7C683ptnF81tb9bd1huNwGikieGn4
YZfgHoIht/GwfsM2bbRWIR8Twp3q1HCMUpZn3XxocWMR3gqu6x0cGrAdf4On52naWROtfs1aU45b
zvfwQ79OcMFp1vp5lIXDOJl24OneOCdMJaU2QkKav1jc18+VM4O116iSYksf4cc1o10IwLmrChj+
wRzLE7OW15msY+bxBKyLp0Ur2ZT1/kX2SLpWVk+k3WX3okdM6LYcEuya3QIqoKD07KramPGdMeN2
xWY0beiSdIbCdBUONcbD7o9gu21J86f2NVU3lzMzbyUk3BvdhOcNwyF1rGpYAb65l5c3B2ZJqu6r
JQf/lJvXzq8oQ6QY4vAwS2yCcWZutKgIL/bgPdkaQ201dm5k9lbjvEBnRWCqAVdRd21noKF7t8X0
qnOEk5i8Mds5lNvra57gzz4x6POpVB0S8prwcSibmEMOX0RcCbVHIBzqy0ZFAfvqQO2iuog1FGEO
xm5NKag8c39JTsieJZDtfWoS7ItQNMfj949JfKLcajXqMl1qN05y7DU5CnzPPC2y4GR4CnV8nk2D
Y2RxVgDrfiNkmInZlPyOiVc1W+BttH3uJ9dokFfIWiRkVljIpRTiPBlo2Wi/tgrG/bEXiyC3KT9x
E0QGp82TvT69rzPZlTMtI4Ei16R4EjfF3oLfiTztfGXs71x/pt8eRWH9Mxu3GNOhCfhw24isdwl/
Nu8sXo3UUYweEbN7IgHTNnbQT9QEsGuMYGcsf759xcPE3Q2Cdt5Ys5tZb4oWi0Zi35HJvAV63j+I
fAOxWILqaKRxiXO2BEh5wSQBK+1/evTqZ/7ju7Y5qeRRGwQEe0m50GVMRVh0r0M90QTb6sjJrqy6
r6wKwElBdS4hr4KE6eQsrjfE+4lew/BhPlk1m9m+gP48eUaiJuHqMPU7lr4az24n75nQKTYjK88r
KkgRjlIUZky3bBflSqbBhxeAyTfC0/msi8XtU2iQGEfZLq8MlA3uS/JHd2zEYUNZQrocQYGLVZVL
Hk1ytSVbIerEoJV5WVGRKLGOsVHY+D75kQb23B9lyhlToYraCjCF4w6et0Be6pbIMc9ya6o3U9Lv
2+mSXr2QLZ6tTktMlGm+40UKyzUQd+HrgsACeSNY+V1w5y58X1a0l9iYS6DPfIBCrmuvAJpYcwmi
slDU4tvKdqU9fTJ4uvaCXIyajm+f5ewoZaWf+oPsYv2tIQY1Wbgd6YjhinyFpj5IdNijAUE1Rqnx
7/ZDDhA19rxjpcrEonaHyCymBdDgNyL3FaHUN7edc80zWBOIqhiH0hRgBpLbKIAuDAHRcks9QCWx
Af7DPzrKQGuu3cQ+jwAx9xLxmvajI1dndAKlNHwWDj4/6hw3jAximy7G8DfnKW+KMpu1LNxtpAS7
srNIsbbVdKxXWeoJLs/RoGX0RQGncEHgWjLAa00VLUzHtMteMwSB35ZI1WD90pGe+YWYNveqjO6M
J6mcx76YKzDDFau5yTvvkU4CxlfU0OMU7625jxi8GBIox1ebds5DdOWu/uGwrdvqktkAY5Ekm4GO
nQtXdYwNyzc5Gj8SaG14+LOvo85SZ4Mm/UWJyBYnkWTE9qHz+DtN4UpVh9p86en9dBOOWvMKExWx
I6vNA+z4nmHXJydb6KZXp3dNtBRh/duB3jCFbzsZAs/GF8icp1QVeJgOmwnSqv892LWKIVAn5lS0
BeFwTqLhRZNnB74lalXBD/3r2Vrv1skuh2Tr2PSU34jlz4dFnMYOgP5V0Z5J9QcJYZ2MTxAs/37v
87gYc/j8zD2Zluz7WRNAv90tdnf8SEiDeqHw7zhjG1qd0IXEKd++tH3EjClxsakmfJNeOE3nQzDh
GZsb98wAohKCA5AlipZOo537bTfT7OUI58DxOExaXpZCC3pCd0W89vY9xunIP/4yHbxTh1xeXcH2
1BXwVK++J+2XbvR1qgZ2LMKAJT/endZqF6IAEwuk35KRsQzqdcWEPDS20TvGR0aRfsbW5ieVS/pl
b9A71zbYe4+9FXyvFpvHsiQe7pxaSAH4BQfttmGQNpwrse19Tfn3NyikKkCfDCORo0kyPAWLwo15
Bx8GLF9JTAAMQoV9Zc0m+b9OOfy2xOQ9NONFTRHKswUUsz2NIfFLpp7+Di72VfgiS1+ZoyIAvS2Y
L82rVkuFgGAUpsz2+n1ndPdO4GCwGcNCRmsrlf7hmeokWLGfcCQcVEqBCIu9fnVskLCD4HiTUzAr
OffINLLwOJ/WWlWXJrWUxMRap7lKhYDGd+m7PloeoGMrC0xPH486T8iDx/Gke1k9jk6TlA+u+ATx
44J+3xNKN4tf2ze4KVHIcMTVfN3ApXSjjqNi/QoPef3g1zUaKgXO9neftz3G7Yd5U2Lk3tj3FqCQ
4eYj1RKT2WOpYv17Mv6GFpaTpt4mWmB0YG6fy/pyOGhhGNbTriZZZxxn36ZAU3sJ9LMl2NDXDe7Z
QS4LtoYbktFpENNW8EMjSDSoOqC7LmXkp4dYwMDtQuLKhpcmULor1qqOT+nq/xACGs6p60C4o+2v
/UhrpPR29yhE8rYR/G4DA7RJMQhAbkeDLcihWzWljarhR1xlYIFCBVgvmO9Do2H3FY2EB/m9vZ8o
kn/TAaMEe3u4Unlv/PcBypb8hUuoA7+L8dqbnbQAoKJIPBTqpeVHfI0kEMICXRQPTwqJF7IvVOHM
BTDE0EKj1smcrd2RDUtWbWBbdTyqB+kdzAf9+eZd868IzbwPiiCgrQvb7wPMoRI6DjEvwBTxVoIW
J506rPoqfKlfU/r+gbpeCxWpP5xIsU7ZyY/4a3C+SRgJZXHy4dgFb2F3RR/joLcCFyycNGOsDBh4
cmbrqDKMIEJsAYzjJak9OKkpL+OWtropYCWGIl1yVZjvO3hnL8I7/6MPJW/ogTCCT7gl1PI6r07P
pWeVPdWKXaNsNEZ5sctE86QAQMIYb5HaKnEEchXcf2Nprz4fa3tbQIG1jrGmX7mTFllKk/WBwSFJ
9529n2JtThwwJw0+oqisw8InLq1G040rg3aeL0Q0VyNoYNNU7lj3VogmV+P8/XhzWdt+xONynTYV
NUjaV4pfWKeFUTp/VtyD7z8qAc60+ZPv1pmSoTCc1wOfcypThHdjzuVsAoJDgd0rE2pSMzygm4Iz
36Mb0TaGSw8cM6i6y6VXdaE0+qrBvAuCOuKdWn6Jk65Yzz2qUjVUReq2N34Cz3PYsjeiI2jNsbmO
xRvH/BHBloPS+2ubhM8dcS8IU0FQEG2DAXl6WpyjUkBOT17FJA/Rl/JjhW0Aoi4XQhfCCkMrbNb0
72E2r+WFPUFwA+wGezGzrwEAnLs7UDFIJdILvuVWDfCjG/acWvQs7DwaNirmYiKmHovCmlDZvYxC
ToKjcptIiPrsA2zCTk9t1TC0KvRoCBGPqCEEwsvoDs/tiHWAqE//i+1lC9iZtW7FqjT1EiLPya4x
mFUyQEJfDT1OuG1UuJU3rGcl7piopMAeSyPY8NMDFwrJcXB7eVq+FnK2B/1716zKzJBsdi22z/c5
AFHE9Tm5N5WiZxgNDIfMmV2YCI047DYNA6qwubUSkAx8R2RY5obBvxZKjN+dyfU8r9vM9MQNe+UI
xmCKjtV1wBBgtO7NYzbXggPGQH6tPya7K3gd9TCrMFBIRQ9r5fdslPqaFmCLXnWm3qLi1uInI32h
CNt7gTwZsDcOspNclBcuLzHihtC+rXAyp3qRhlTBmEbcEi3eHSiTmg9jv/ahoLjDuf23T2/Cv7IF
Cy2BTLzGJR03iRL4Bly+kzwjYyrILTO+C9NlUNMO7hENRb2t8hoMj7iBbnPDj+fxdsZhTSGCd+gj
sgDinZZHQlNhSp8pQQ3sVqqMz68Eu79OuKJrc5/DTx/eZNUUWT0dvs+clEDYYMhxDNV/c8461qSZ
rENuqKiFZTbZ5iubOA6FYdrCSH2TbNNYlMTIvfC9h+IG4lSDVs4VfOjbj2zDfFVDu6uRKpHKj3ZE
0+oREvUIPEcJgF6XnbrmOVyTu4oGdZcubuRhovVPkMYAbX0shp/IrpsUNkXAhfI2mDnUWmx5Jk/B
H2BCMo9ZjA9e38pA5jCQlT9ujD8Q+8kln9DORtPQmzGJY/9y+DN93tpY4knkeQjSbDG1caggSUn+
S30piQQhoxs84bK6ZKPywuQ8p9xaNumS079dlrj/hykFColMbCuZ4x37yDtZ/Rdw3hD4ZFDIV5FH
kA+OmGVfEZ6T99MCa7VnwuNVKjAD3xBNxtpnRFo0+ufrsH/S3ua2EAe1HVrry2+Mx/JyZzlUkfdm
Nyp+RSUvw7NykQMQ4e/6AIZ9Oav/G05ANIptOvM4XDqkjyjZhOsegTR57IuM5CIM7St5DG6LT97M
6FsVWyIT6EaPrwaPwwsjqjoawSHN7Lx082CqobHYli804ecAISoBNinz5S06OH1fFqI0uJnQHv5G
KCvU8gmyNWXfarK/06xFme/iIY6RNalPrGAzk0GhA9Fh0xrv3Y0gcKyYgbsi2dx0XXTvc0gzvPQp
ynVwenQWVFwYigAhV0KxCGnJ6lvf+guunrlJ1S0x++UgTgtNLEXdXs8V+KQLdpHiGC16kM6OqWBc
7Fxmf7CRZtc+YJBrl7wmsjh4W16cZOBNARC4x4rsCNsknwgdx4CKDc+MHWk1wQbD68PhJ32e3/tj
Vd6JhCXgUGEbrLvGPlxC4HP7C1Rnj8P1GKJhwFvtEcUO8Cfnuf/IlXl+se8N9Bd5XXNzVDGM2YZc
DqIjfdBw7AFEsJ7Go/wtHBuGe2+MXjYPkZuWNItrlWw0oAvpYMyjbonrS/M86Zlr2qyqJbceFz5R
h5cNE/w/uaGAQIV4rRBN9R+PXQ+h6et00UzN/LP113gRMy7aFN26amj5xzMt38mIQfHU9IjnbgCm
yfg2kRorwiWa4lB9YGUOLpMsuFtHsqZXgtS5wt1CBDYg92DaNUwNkVbVCZhf/ZfQ+++ne26KzWDP
uOtmM6lntXVEChz/dUo9TATww152ZDtJO7904FNNTL32cQJ2SIaj5Q4basqNS52Scwknl/fsRyBr
B4py/G4z0SJNOC4ZVKnvxn8bCAfLbC6ui/vHFvUDFm2U3U2MdV0kY52VmZcg3Pky78zG+YiF2mI3
9DbeGOOz5pdNiyAsZ7A/cfgwOG2OIm6R31PpJGNAu4kTAgNBFpqqAm9IXwGHA4JnbaOBDO534oIZ
mPZtH46/aqtiH7lJZKAxu0M6x3uMQZ7/0lYalDfUZkij40LGqrEN850BO+h6uFHzcZJlPT4Q5vOk
6aNmDvTFZoMpQ/fRdAdkyPTuASpcjSNt+nrOHDbbDqOtu1Hj/eq+nZ7uCK8ku94qLXjAvhNlEjf2
LCEMQcCMhuQLPvD180V/2DbxSsWy1EgrGth+8y15gywRmfNicPciQ/JEB9Xw1m3uAH/twTDnothR
YSe0e1oDp5miv92ph7XmBEXFFE86hIj0jOSXTLMzi08DWDEGam26BMCoe6sYWhqA3Se5N+Z0ak+a
hSUHRUqrtg6dOHX2rHJe6psnon8elhzwWVZHZVbB7p00PjLbgFTeooSKHM3IbryZ3mGn0RRotk5N
tciGk05xzLLWs9cKauoUx2aGQ7ZQ7dDjdQ5Um78Oza0AB7Hlwsf6hERwmB++rCLOT1/qv9Uk1YyI
xIo7vNHVxjMwInUCnW4NKrkB24Q8J2VnZZj6cP9C9I6J1auC1ZSgMcfHnjINu6DGElG4PIOrWSMK
f3SpK/tHR0NKYPA7rXuumAAIwRcYVS7kzuYMLwgo4+k7ZOKST/kCLa5MnbshJkIBK9Ek4qon49uM
pStleIZ+6qzZBkBmqjJfMj3bLRBFkBM6HbAbqsF8m+Efe/aULKW1MeZSk3RyYj/+zcO8OKjDlLmF
o/7PKe26k3vj7ZZDCXyuo6TyXuuK3FRHW+M7FG0t4Qrh8Wzn+H9FZ0XoWY/oKW1yx1FqgrAAbLAu
8ZzniI1K2J/BHbPaU268lO109RY6ala/bk1w8eDf6RewvP3qK47ox4ydFSXpI/1FHxC/N8vcLvQS
gd/LZ1DBYMxYZOC1QpVCkoPOWO+bQz68mgUcwU69u74rd6VJYBRrwYUt94jkTf2uwqd9iBXY9W7F
wFnoLEitZQyjP0YsTobq7JFlJ5gZV9Hw5ASq5PSlAqA8YQrS3/fghgAhlMPt+qNH+q2ZQCQTxoBT
8oVy1h0ic+1m3D4Z1KhJRJGq7BxXXbTlszkp0orYsu/kgoM18x9XcKT8PO519loai6IHkeFfgDkp
L+s0IBPYbjpmB9Opz5evePIyzkbmq6phaWVkS+YISznlYe22iiixdXZCMmj/5ZRTD94jGWabEG1R
Z8FpTpGDpB8E75DdmbTxiHIxe63zQpTXWcDPCFNGSEL7UQLIvZ0udykdzSw2pyfBqqgt/VIy7/2S
/QP/mYAggZk1kfMh4MRxgRwh5Ze2CExeLsBw4FbXCssxHVtTGgoSpOsM4U8eFtAI4LaIenTybIN+
VcktCi/q7bsa1UEv4iFfwzJA07GfTtryLWmz+CoTuDP5dUJ0OH+ndGqN1JpMkBX5VAAtmTlf6+rY
sx9hCg+PJ3TyseXseA5Yc3+8YmghRSb6o2/NKaVOv2vAC+m7KOPGG5IyIgsCHKsMbik6QBX8YpF9
byV9uYbBbOYkqkscMYPhcNJ4ZnDN9Aq4Fg+VMPQpgtz/vIIhwi7tmxRLvaKTkA1Hti+wkSLnkjCO
N39K8nAEGNDVPK+C8n1nDqRMgHLSkbrhdX/MYNx6JLUD6tqwQxmmvqpfARzJ7JFY23J0rTLtBlaL
qFNm7q5azGSLYJcWc9cFTeilSwFdGAepM2O/wT6/N2nSGHiGvgXQPqsiRBUsJ7oQXXuz/peD9BRS
vRLBfGG4M82ITHKNIkpe8hWybstvfF9MnYG/i3RDzx/1z6y7KSYCk0n2gGaY/mktOzuWb/gAtoQK
xQpyvoghTAwElTavHtire9Fkj/lGwAl3tTOdYifKTGYwg8qE2fiD7WTDHgzGQSYl3FnU2mPwPDbR
Axsw7a/BdcvKT9WJyvw5UQxws3xuYf6A4uIyJFf//a/mdj+jXE8ZrOlhNGJwLRj84lYhJ/gQIldz
GZp2w7+pjtzREmAIvSYB0tL62UlAStteySHMtQLsWApFbHsO7kPkaCHES3KRscdqV//5gkNWQQyI
YOkFVcBu5GxuOI3Th/8dKYFy028Lh4D7jgEm3yzdpPP7qfWjnQdQsSMtbnqYtowJZi6OWpObEzGI
PsTvuBAFyf2eHu2EQ7mmoR4/AfcOOmJaamzgmdKSnv0c63gSTKi443PIl4nScd0/pRWqWES1RHdt
HB1OEK7sZdtcMh5ItH3QL04iMXFF1nnVAPLN2O7l00nw6bG53LEdN/0GSBbc4kpKf7LXoNvWBWYa
t1zmDmfdkGuiYrHdVkexcLs6g1JdnOvPZsTSuM6dZWQf/NWEiojxGIiLiHU0cReb5eJ7/lT+/7n/
VFlcP08018t+Ce2pd0bTBuIqahASWqEX19XnEAwExhLl+xvMKUo4s0YHNJhl5HdhJiO+S8gM0eGI
+1/CRg/LIfT4bN0OjPX5vvEf0dnURUU1BN/UCGdEHOzYQ55sy4ym8fZfxQb7gS/GmYgbN3Tj5zfd
oASNUcI1vOIColpj3iyiDwa0nSOtm5sgT46wG4320sXqU/vtAjKxVnHqV0o46icS077udGp9C366
/qeU6hA7Uao/Uh9unNYmfj1mg/rZ7iE9QykO94BrxJTH6UvmXm/QTtGU7wx4eZlBW2WD9px7TFyK
Ry/CqqMM0FVSc1QbpOUZXQggVI0FhtAcGr8Git1aaHPmU47MPLn9tIVCjEzWaAKRBhotr4XlhQdt
oA2pptp06mBnnEU4kULO0jaO2CG45pzokNy41hpLHUS5TRnRiUXFgf3Xh8h0hNvAf5RihC8bX/LX
oE/leELK1/0owRJEr4cApquYo+qSlgY3cfdGduOpn8eQZDrzL9JifNlr2lDYb7ID4QOEjzOJJamS
pLVzxl0MJlmPvVvRgTqKdrIrtZO50Up3m4JsVe20zl7QZEooKabWsu6yZ3vFXsPPOs3METeK1TnL
6QjTEV1b6xa+hz0G/1jLW3BTnxtUjwaYswiq75TcnD0j5pwy6+VpQQ7ZZr0kaZ8UmoZ1D6d0MPzz
qmIWDqDxjU0R57VmlLxCoOMeBB/oHdjBu1I8eSAwIZSHPg/jE8XeooNn+um0C+DIodW/rjKzxZWI
M3eVxAVK/dHwpXukc3GS6Et/BMBT7YOv+ZQe/KQXZdesZ1C9rX6+9URpPSDfuLSDhEaKG4eBfEx/
cs4BGXlQMrpI6CmKYTt+HsktDACtnfnOjsymM5w0wfLheiofBHGEVynzphRvtYTu0BGcXJl1vzeV
UR1TfB0ZpLWIEz4nO3C2+hxfhGI6QzkNYb5iBeeo7ZA+PGnSSMNu2xiLLpxslc15oTPHc851fnTn
qiQaYvWhYvof8gAic8oudxbKSlomvI+XT+rCRIZSuFBzUJ5tbwtStEn0zrVhjJZa4HSip/+LX493
hk0s4jnG2e2VJ0c8bRVN1x8bhTZ8tkkJWN6VYW31H49RsncSZju6U5jbfhyp8VW4II+zC26uYGkg
OBSI9FZNk+Hu/7RCVxxUi9pPXHZS7SfgDwaasJCW5NpHrJxMvR8z0LZlQqD6MUAcXgyVh0uHOh6p
jYkpAmcj63QUT21ifhs03IEWk42IrU3J6t4otu8JWaDjNLxKlOM5LE/gm+upaAhSYTk8pEnp6xto
Mwl8FO41nFjX75wOf55TPPWGUzgIpx+71WdPYEoyAdMESTtwU5HX7XVa4vitmF4d2TeUNG4InQ00
5Fio4gVpnyzQhDY1eW+BzOb4wxs/ce9tkJyrucQasvRogky+E75u40483aro5L1ncb3/t3mhNjOx
rMES2KY0ScMzbQGdABiuxRFauLyFElPwdwebD/4uJgSK7TAnrEA22VNiDu5+hN599CRJGRsShpJ0
diTBYQISAydiYApaxvpTr8TYa4/Ly16IXo4ydrIWjIMq4F5x//4nA134O6lH9YNUzVFB4t8rOvVb
CHN/HrzSeLqbk4SfzcIiOS+fLp/0El9anQIm3PB6NJt1fagXiBS+qEWvMBXIzq/SSHZnS0VcrrEy
wVSJt43RWPqcGDHz3n2/l9SmleQdqZBpsrymK5ERNB2+qMPXOJrymmDflby9bH4PqsrhQhmmssKF
OU9wAXyr4/4ZWyHJTQ3xlpMUcQvfvrX6uMKCBCXSxE8O+AUHuRAvxHOYP6M4YrjYeB19FpFXJLf6
vzwVd37k/IYoQc9C8VcjNYO9oua6KYE82JTm6RFT1IIch++TG4loou7i3Z6ho5/ykwJ47/scR71r
B4V9KBvd00/uH/MtG3GGhgM9NaT8xf7cT/Syrx6ftbBf8dZpcSh1Ec9jpHRbfH8eChU8kp23L6b3
vE6ivULgey13vS9csNrMSw7Vdc9vqfKHBw3r5BsfGJEbJJtsKpsMAIjM+859eCw3INLrpKD92AKr
+7ospsS137vp7jGeqNfKt2OscOM4yjmCDwIZ/wazSx//QXG7ebs0BcC1UP6k27Zc01S7YSr9aPj2
cMRFWgakAlceVWiNiK3Ql8WxIyYCBOuaXfvq0VgdsguIzeQirGL6/uDdnwHjTlv3cNcvRNRt27+i
rEolLWHSfOnuwTOHbeCiRiIhoByb/Q/WjU8CxxmbRWGy/VAcvXiQpccUCuMfYtxu9Wx3Von9GV+Z
O0hD+65M03nkmjUjJJSdzaZ9PacO8o0bvq2VLAwsUnG2eO5gMENMRfNxksqOMsfNgv6QJcrCPmk3
6Q7Q6Iw4d2XUuYilgqYntZow/pJ8l77KCE7/drqMrhAGavEMi2BWreGv98fDqE7R0inhkPha2Iev
lJ9XZY7Fg3EGXjr66Gj0+aFVg9Oar27jLBuObE0ShEq7ch+AIJQNFiMsvD3G52osl7eYJIZCrT9k
f7XhquAhG8U8uqMULKY6+0/u25ynqkjb6a8gYufAqjtGYOg98ygVQNKuMzqC4hpurn1OXSYtRH/X
KJsZJg5mI0NX/im70oZfMKLiDpzpt+GvF1Khc657PSrGR5oDDn5hiTSpNbbgn+PVzWnAQYKyenqO
L+O4RPDklNgyCLrL7YFD7s/3q/0v57JwCyNeFztq9/EAWDIZkvBE+y4xICL4MsD/ZLdgqwCHYvmt
q4+EI5OfPfkh+OwaclhYxVzXTpyROcMXXYnfgjDJmrPmsD1TuY2sVLlElRFZ+HPQscqC3AX9kups
mVYaQPDzbJk8K9wgtgAKrn4PEXXmR46pV1sUGc+qXW1Q+MVtJAVx4zOXWR6l/t41rJH2JwSVHdlp
Ow42jY4gs96wbqmi8ESAtCsiF7EKU4LMfwn2A2pQzjdYtqUagAJv7ubiQOkNKrWKmkCVNuHl+UJ0
Br3MahmQBGR4aNgyC+ROnTp7Y2ohaV629e7PfVF8SLS5pjJzVMmvwPhMfHx4yoTq6A3ONymdPQIH
I1gBKqlEDkGzEiW6RLSFA4QfuMYAEDzgfXNexJI4UYv3oJq59eZq7nk0jucqPpkrba/zc5VS+XSc
Slj0qirjeb88tomOVldZQ1lm3XBh32tRt5azOzDkDKwnTkr3CAF6kxWpkyxBe2L97MXFxbeG7bU0
ApKlbA1rG0OhuPaTxYl75SEsUVFxjXRQLBiM4OLHjIfxCG57nK2P7WKEeXI+z0pZtJjSZDWde7Lr
DO6nzQBNAekz3j9E9EwvtkIAIaMYeGMCbBN8WVeOE5t3cKikh3M8mjyL6EpQ+oZfqKM7gyy5o2Op
KQUt5PuF6sSOneFE8iOk1WPFbz5dZeiqYBMWyLvJncXVfgSK32PZgpd3SwdlWNdSmerpTCnpvLdv
sMbIyiatm53Gwwncm172PY6WVBvi3dI7V7vRGfgvoHoL243nSgAutkS+JDDtYHn+sV5+DxVOen6n
VZETk/6ctogJCriG+tuNJmdMMKN+XD4uiQl0wqR+Uq3HjeDGLFUaXaHkviIneXHgOfX4gsAMOnAl
kdIti0OLWbY9ZAwLWH6Zr8+LUkPPSzVo4r7RECMA6lrubmr7p+pvJTFq3orOJolB9ZuTF+626Nga
nYMMICilfowVvwCfJ3TobDOYyrO1RWfVxO001eKiwQg1XUYGFf7uXmvp8HzRatJCScz4jhXeDW/3
kMXgdhqkuDygBLvX3Zr3dEBgdxJLgF4LlFtozeyJOL6TiA6e8Fre+cPSbsmU63gibbw1W/7lzcY8
to3b5qbs+E93lEKGDYLjawTF3I1Rtg3mNVvulVD8u2h/0K0eRIZ+YCq39ZPR8iOqRxtij9WoUGFO
34RKsjZ5ZZ+Rn9QuIzuhoKc2ybAG+qQLRhJuipdNCV77ct+oF8NltucyPS/A9urpaMfvI3ayP51Z
h19ZDeMqSdGUVajgj54SKKhk8Bkv5DWVOhMdiKAMF2kbjlQdDlr4lmFdPISRRrhOtwBD5LIWVF/a
SjtxStjEu5LXDUrChGiFh1DODTC5uN7BPNr7WAq8Rnltk6qPtxEVQAtPRUpwdv4WIdU2JGehlvFN
LLQAncRJ7AC9ix6tsjn5w5BP1gRqWyHxDdEGLLPwL8bf11wljkPanBG/NNJS21Z03cA8OByg6UbB
af5sT50r7dk9Ulf7wG3VAcFJx4zeG766A1Pfrsevu2guWc8LtJbM0r6IuIuZFft46gzHH9UjZrJk
rRKJt2iEXEt6qFIBVxZmA80Vmz3CTobyJPEsvUj9OYmn6ju/V/Z+4AE66qs2ZVlSyqps45i0dYv0
rBQu3thfy9wwQ6GmXrIKeoKIr0QhNvQQjg8v3o46J5MQZxJT2jPU8xEGVM40NH87XjAlkdNo5luf
WFgOXkKSOdmip8AaGJ2P45vKyrCJBpBUbK25+OvKDtfAplgJx3xRm9ny9kjmV0MnoOF+xLh5ggnI
1QOwPqGU49kS0I49pWdRti7M4GTggXkYLfGo8uUFZcW/j2l6okH1kztoktre3rWwSHUqayui5Ai1
kY22RfJdThmm4qm4pPpOO9eXARqN60p/nxAir2zxXo3fsBYX3CYb8FH/R47qxU3FJZHBOrPRrMfy
/UBetjG9W5dE7fGOpt68xz7sGBqhFU7qnUO5KlriMkA8rJq5mB0Vfrd42Yn3uYG8qRyNhkoqLH0M
2wR/i1qyioNXgf8PwOJQop2v7Wx8SevML1ml+U9DgRQB3TyY1A0wAtoJpZ/zG1ouLAjzhcDpHIWi
jjxUbyzvH5Fmg/gb6jTJo29wzRwg2uITLAAR9BsyTHbYgLmz91X4GlRF/I0k18QZ9WBLmxFyFpm2
iUR0Ynk8bZNDGWg917Cqhmjx9oTgKL7d/ZlkpXiZ5N7/zdhdeQZwVDKSpiMxanpP2jziJLzDs3lM
AXR6wS8J7v/WWrU5Wku44hT1jJ/vqF7JjYuxFlOn+N/zwvlqUUrwyBUV2V/w9tkiX6NOvn+am4rh
tfnKoXrHLVlkw2S64L7vNGMZLNb02cruGpG86XbS5P1jQivp1GqTF614dmN62bplCPYQ/PoiGp4x
UDffS7CBEy4Nx/58yr3gmiiWQi/tKZNK4MO4ITgHK1fUrSGlAn9LGHcC+o6KFTqMZoUP2PtEGTbK
9OQmNCwC/2VzEcU+QpYZ9ljNXwYJPBJPyIuNFn4uFeK1uxfSQpytD6awO6y8rukFOhgAGmmSB6t0
oMQd5o3Il+suUPvPebHDoZJVukQejkuHauswX2y32VOI2KnpmKJKXIxpNmyGoKNX7tCgv/mGakEd
GI54qcUBYg7EU4Z9at6bS1vZD4P7KFMobcU7ZrXlFlna9w9C/AfPVFDbaMheqNhCqCIQTO9lbJm4
lOcC75LtimHRxb/01l79dAAiPt8gnO+L6/XbJJFipKKockmZiiV+gnZ2+/e5J4K+oGXL6sVoqxF8
8+QUXaG4YIur2rh+ePmSZJvn2oTwV/0qoQO7N3d+o3QazsXPw1mvxE9SNV4u1C9cqzMHZiVyX5ce
d0v7+tsAT0DtRNQE941lG4THFVTTsYZq3Zh8vbupjM/dSmluR8l8f2uH9qS5f7VJdyEPto0sBoV/
iejceLqN1JzG3W8UFoe+/Gu+l5MCCOTAcKO9AEpN59WlsBr9jUZw156eTorGRVUpbEfKK4cSkD/a
ZyndJGsrrvFANmVcANeAZisQkIlNYu0/QA91XxVtwFbqvmYdBYCta2KlLrogfLom0rbU3gtVHOUq
akWZTYRczfgBYjXJCzvu7VrZr1EcVRHJ7pd4LcMn4IMYMxPwzxtQfqpWmxuO/+kACttn1YHqmhVN
mhPTeAIwz/THXWnSTwynMbTTGn8AgAOA/kY7s0JMbaNE/t6R2NLX131uDj30N4MqZW3le5q1Te0T
OeHzCSTi/7ioEF8V3tferEhSDo8vmCwe9Z+HVp+LlIWn2uMjj94sNoChEj9qo6jd/gSvsmuWaaxW
CmOfWweE+p1lFhIy4w+I8nN870T1jlu8vk38bQD9+fao/OGYPdNuhiiSRaInkrl0zPsKccOJSeCm
uOQ+8oQd0h66nTxZkI0LvPXO/aW+bhwMLht/97BUIGIrvroimosoSfRZJ9SS4RfuE889C3IO+Dbx
uDOXd2ul4o7G7qF0JizBqRvznmY2I4+kzjlqVAAGCCe/2gZvFsUm6LJq/+lxp95gnf/iR7pWjuUB
xPiWdROHlgRE4+4yw7quiM+PXASgldADXnBLYjfmXZoZuip2Szm7kYAhtyWdwueBa/x7u8IRNx0i
GD3/CLiPna2AcScE8xjzT6pAI5gdw4Xcq0LlWL7txixcjQF5ndTzNV3l1/VWp5Ys6q66lnvhmYVs
ajP+8boOosM1gHgCzzVet9Xc+V/Da8r052qsNraxavGEAQcWXiivapWHpPV8u2x3EqFrGxR/WJA/
yOPqhw+y6JXg3sVy6RGsI8R/nSwokCKJOv01nWbNtbYKnjxG1rJuEBZjWSmNUmPm9ZKgSptlyFM7
jSt4dRCuS8tjrDX4CKwQal/q+j5UuRxpoplwNYQF3UK2L8IH1zz1X8U+2H2BXBj2Gsir052HRNAe
6WRtLcJeqymETdwPubQfFLU6yYMYqYaEZ3f4raLvoEQU5F98PxlYr8h/SwXtp4Cwl0QuFTHiRIHi
HgO4//RJF5YgJ283QiiP1g0+5QNbAyIJjJzdc6LjCKLsXd0MTXIbneBG4/W+2Eib7SbdLL1eTpvt
AQOzUgnIEkGSCnWpmqCg2xwFHEmDfYy99oRkHp80FYCnrek76SUSWUs96NFCp0DrzRzxCTqktmix
z6uuqsieFx4cf/yyOrKTRuyzMMYV8IB8TzewT3uhqwYOAWgpbJK53+QT6XWvZfPvg6WsdA743Pyy
UjDzZyfIxfAz6Oo4eiN6/ucP9D9iUiwfDuEZNfSMbtf7q+3aclIkhTPnYq1v5mrKino8UJfEI/V5
C6yjyl9ZfSVKy5pDDQkhHyCaUlHcaCbHIIju2kQasgCbS0YszjZFGNf3WtMFyQeep0Nl4+QZAwas
xEKLEDz4ISwq1lN61+YSCP0E4rDZ47T8X5biOsleBXoiqtosA0hadu49i1eXfP9Hkz8BUYF5WnV8
aykr0S6aWQmTmOjGBWIjQ919xtQ35FEmdOfuRfHn8guUfWME7/2+7dc6I0DzS6/9l2ifC9uyZZBw
RdHqT+cvQBtHNG/NmTzbe8fMCcKfrDK8kosdFYPjUGUVECtDttnLu3diZyUZM2/N3LTg6Wg3tMTw
/kJ0ipe2CEl1WcDU6pIk95jGVRbvSzJ3s1Zdbet8wKqYiwYfgETjaJtErph8cRSGzSI9FTE8EdU7
dwSvVBm10IqXc8vVPSK9XBhEzlnItppCnEh5vIoDOl3dBkpChwgR3X9XjTpwPvtQyRzmgDU5z97y
Z2q9iQ87/cNwPnPuA9IwLSy7eBPln/NEA/nqqM4jHqEF2rdgXp33VfP8iCoXiKcSVUPYDp5chcrB
DJSM/BBv+mH6WhJC0s16dp+rZ5xX2LonUxXbIpIeN7FVSCI4hhMrNozRKensng1XdxWNt0uJyWxq
DKPNOFq5ziksoSJ/p4tp46wtfUywUXpkFCGc8DUs5NurRD1wKwwZaZKjeAYTs2RqG7tGLUh3xjai
kNpHlDgtl2yD5klDyX7YcagNiFzyd4QmVMBi/imHeGpsZwf2NZ7kmCGCn/jB8AqTpzm2Mks4Q2iP
BpG70oa02G9zXg2yDHY0wKZpxiP8S43L7A08h38poMIXcgKDAx+DgB767Xj0wgK7rvJ7S3aZ/yHK
SWNAY2VTc7dhPsvrQ1vDQTlm0A6XG/rOrxZgkArSAMlLhDNGeZL2b7wdWpZvHGxRnM6k/ZT7t2+A
LB85YCna4NO38vNMuAy58F9/5r8cDi7AK4Y2TZgrcy3cZ/DqXG67awA7pfseGMMMJDx14dunARIv
brstRyOZlJLmJ4XbMZpTkPJcSGRewi086pCL55DE4DakO7FLKJ3HMqD/T9wmWpyqu6EYe17H+iSY
spZfbqThdrOAwF7k+qL0QPVIZ6Njhtr/5Mzk107s0JKbuURg45UMLZb+2y37AS++IBum+rMfKZLu
Oq98g/FDqkrfyVv0C4wHqe/Exlbzly7cGxOxfdQnjs/JWYW49GESLHFTIuXjctJD7RLGsRtZp8JP
pV58gFPjseTtXwql0SzcYVD5xTbJYgBvxP979v0VpRgN6Jb+KuMXcYas8Gess9Mg3rWdvP+3kILo
1bO42LushOVG+DPleDYAFKPhPFAreqY4RI5Zq3a3so6gh2o/rE75xez6sSufBXGe7Tsk3qq7fkO1
Gz7lE++6m8bRhmOcUrtF/RWwaEVGjt33Cd7dkcCOUW7tg3geW2j8a4g/ztEkAmiHr4nsFvpTDtGC
MyTWpygZw/SMgVuZTXt793mbyCII81OF1o5z1Yvo+VcOtTgTgrfcuyElO/8RzOtX7UbqEBrNJTQU
XgMMuvIG3WSxYqSw/3nZYd54iVPOZ+EthC3iVRJ3ZlA0MUayq5pGjFSVEBTTiTnNy5rsjrCnxvQL
NJ+flNwDpbeZMOzU1yMVhcUz3CzcbbTKmfwIPvW8CbN22ojuWhpap8sl7Dw5a98fnGV9s6Ti/Lb5
7XfDlS6AFtrJ8we2xFqVSswnOCFKzTFAkeA9W6gIhn4zA9hJWjuiWv9dXHwUftZlTTUNoPbVX2/U
BXTY0MYQjQCuCEDgNhzLR7a289cquhM5h1WjqMnuDBCLXfTgWUBz3k2Rz1XoI3bJze0tJSMGmHYE
INgmqIh5ESda7+LdlFRvVRM/rW/faj+u8ocqB8lDiirvfmOVgv6Tp1fT0Kq9nTvUtAfBRi2xHgiK
WeIvNmkhCEFBrfNicefNQBXqvv0tthVW1WtRxSU+LUA7M1OmULonz6EPRpiarXsbPZCBfGElJNZJ
wi3FbsZhVtPs1MTCO8Nva2euzc8YSi+5ugovHgfs+JImEXThrE/HzIBJqp1TkPNNdf17W8hMOF+Q
WFUeoINKju2TurD2Yc5HqSU5ezU+mJI/c+POWO8BvcpneT0ivI7Z8Rbl4MZFFNTBQQYhjZbC5y6/
sHQKFk5/SeBhUQeDf3vtQw/DcQBIPhM8qlsMjKMBw5+SLZOmWGEjyiszYIuK1igFzchq3r68IrTO
Ot1rHQQQpt6xHnW6O5calgC6eqkLENeClD8wGAWhqo1STqRNDz9RvH9j/UWVMPW5HRHBQAkwRj39
BH64tPo2MorEse9IkFRN18JB1bOrsjDGOa0UNtqTNDCiZaL19v/ZtxwrNWzvO+aCWqB0T6WkFDwc
Z8R8hC331M+qRe1S1fmkd/dDEGSHfVou89LYL9xgM2rdXkVwZzKhbcOvUfHorE0NK19SFe3UQBP8
uNfSPKk2DcA2ij/+H085Paj/fWEHgAgMNKRCAgA4V6s6tXcNNWIHvWF7miZ9656LXNh3fqughWBP
h5RC+NxUQBIjkdt5+gFhOrPlZezBC9NygDoX0rbFrKkEeJ6zQWVM1Rwn4CIhWmJuIkFkHuhvpSCj
ZGUGatPSXhTi8EcwhdxpA0B60JiBk4qKeCiHQo0VEq7/Oq64FyUD+ebGPe3HlhrF0/mvedujya3v
IvG1jLPTugq4TZtHjVUohN4jrCotUxCCgnwciW5lA15FRtaqYRxB/2IersGdSCr3NtA39x0Yni/U
fCwRGIl58iZpCwDVDz38xB+TTuHI70neGV/c+lwaECOunPJJ/jqF38JcUIOVX75uLvCjdCkjUaYF
4zSMavmb8ghjBVq74lPQOgbFmmaf7yfqEl6EcjXbEs5FTyJ2OzhXV/i0BrNl3Vr5JEmxvgdFo98Q
1hcX+kcZ0QiMQFR0mpPlWgEE4ScNtXfKuUtw+ifTR1USzdQytfP1Y/uooUO1T7uyRDxQZqcVZoAf
SfzTTabE5rQzxcMTDGcvhcf2ggFqR8Rbtl4TQtboDuD3pW4ZArKZsQqCQLOpGC/oUJQCsUCLhAuY
TOsmi18wR5pw/ui6SKRGTDBDaHgIKujj2xI7AQQhqEVrJ6+ZPzNjdErZCIMrd3RJsKh/F/8ckj8G
PkltWlc+Xwxao+5WZKsxRac33eEcatR0tdFc29DLmAXMp7U1Off+9cH9v/NfSMQfF4vkxdO6MPW1
/fyNrN93z9Gnr16UPlLfmlJmlT3Xx8vOWdHKrx9v4Pvg49mouzrf/11WFuVLzgHNiX/jhX5OiJKz
07z4SaKdBnKy+GCAzIbTQimatepBTXClEiZF37fMUwuyw/HLXBDmUemQ2WRn1guUgDRQgYgJ8sXP
6HCPzRTj/6fWsP5jTHQKppizC1irUANO8xGRARGPS2nYO1LauHJm/qPYiR0N2/eOlVp8zYqvzNwJ
SCj1q3B776XQPmlCIEbUg5jTPVuenKGVQrR/pPbUAWnB+p5NgaXjTHbhDHr+k0OrflCVOLYt08Fq
khbmAvkSsSi3HHxHi3iIOkDybVY2H7dlbEQ6IFgHOdA+0HSrHB5Pdnocs0bNA5KTA4raohnwEir+
Y5b3MxU6mwTfT+SzaULWxzjfpgK6lceHZTE9GN31cQKrWKGPkDx0NdMWCM9Ly7Ioe1FNEfyYIWyU
rEPRPWK0OcDiSl3qaAoFPHPguQV4HzfNHz4d+JWaDdR0B3Q/JYrOvh12t0B2UvB4hsLv0raCoVGU
AAHC/4MHPpDWkwqR6UxlkQFvJWYj2FUbaSMkjZtDtlPjJr2AlKdtybIq09IWyEDFUbEtG1dsj0oV
16iunYR3oD+wj+SMbcWBoZbOg3/vACJ+stcjKJmsugJjtXV2MkgPGFaQAU/x1PIsySzV29eB9itD
HCtiwLOgRh0q75QmsCvIWfgwpzQtTX1x/lGiK35gixkp62m5f+7FXs22u5q++kNQHuDZWJj4L4ZI
wAiBWkI9UJDj0P5PpOzECKuaeyUpcWuwzjriAp+cwMrEzG8SkRljcH+lK2OgaxU2Y9IhizRcfWiX
UvBI/6Iw74jy6UYDGTxIB1N11ZeRpMNY64tCQtLIWDjEVi/xWbXrnfvGeEuMlG/LdKc77NS7gEGv
0DiXuorq2B1fAP8NHDTxCyLHrHk15KZZIdVPiF/ak7iMMB4tYAeQrmBAIOCd7gh4ML+bD/EyxP4Z
pftEMkd3Xb9eqIsv1ekTD6XmrZUhlBDOHhHpmrMIrioLaTq5cIcTvi54tpAj2JKPkfBbqYueWbcL
o4kj8LG7TU2Igrz2FKDIjUQ1ttuyEOcjAAtz8xupjyL8eLUO66Pmcd1ZujUQcLfvkJc6hEEEvekw
oPe9L0vP/wp5UzAuuY0HsTxhhC68RvxdjkLXAVuWcGd+MFDWryaWVBaIC1guh2ybdw33IJRfHYcD
b0zuw21dtG8BkAXAWg35jqG3rVHxj7J3Z8muoHBH9uQQGr+ndRVmM2ukuH4NDE0gCtG7iIchXaU2
00pkJzLUXXNtu8F2NyAqD6hT1QDWsqi2EIMF14YccpkbUDMPebaGNPehTZVY8IT81zct/hoBkKPq
dhMXnoaY52SAKrX9H2NCpVX/gAZ1gz9s3Lf1IDGy6MplCsA0bzhsr/sVlfWay5922HQcc8Y2PBiM
NZ0wb+fRC91ZCE278kY5nxlvXrwR7GTwhAHt7cZ/3gBhtrSuyLLyLFYQbnSrSy00gxnrE/+A6AUW
Sts3QrD4E8Agn8rdupum9SY9xfzVec+gyhgfuDRwyyjRzgTMEeauEAP4AxXBaW1keIeKyFRMnnxi
zxzAJPJCf40xVNq5h9jL/hIfmxQdlnJtNdkj/nXJUej6ZQfiCkefGJcuuCmO1Xvs6FWk+zZnPPME
qhwdP5VaQbfDAuIx1x6fFl0IHVlo3v7kYp6bcgjE1Yeqytth2UvqagKoKeyaYdHEQ3KPzmP8cuvB
aIR+DOhCbK26CIqIajyWp32mevXKJ/6/JHT8TqJBUfl/hckOkNbssnkjgFW+T6MKhgh7GTJyoIaJ
fAKnkRoK8hmyCYA3g/UpJHtvfL4/mXHZI/Rtel/CMQePIyZteDGi8JD9R8e7xtAbSXSVMZ0JvuSX
daG8tB5iBcyA+CPJgh+OQtqdwMC32xSOFkRlreSE/Q4pQgSii4cAhONk8Yl3R6iUhiJ0OqVGgbX4
dnmm7o25FTqhN5c2y5ZkFPFBW8eZwDruizo4L1uUzsCl4ciArcz1g1UvbDkPDcVSbacJKJwOL3Zl
3cdeX8zq/i/M7/Eqt1MKICWR5OEF6dtziSxWcpzeZPE5forHWZgY8aGazIhPh+d+K+qg4FwRTNol
iDD/ngQB5Y2OoQU/pN99NlcNFcM5LX079Z1L0n7FAgYkJgJtQgukZyJ2TUPLfPl2/a761ERfC8RA
W7R/1S8I3QE4Xp5S2lZEGWnqYlaRpOIsSWTzCSaZQ6G1kRvVWBosAN7l8D0ncoV30VWo4BaWOyaq
WiQ0n1L9b1Hwo3MMOOLUBXfghzDiFjoAtlP39N36sxcrO6jMmxljUMBYlxKx9ijO4vWDjHJUgc5I
hUIAL0UIcLPIFY030kFKZg0i0kLXZ/5MfsSNVdDr/Sng1WWQ0oS5ZG+U6ys/5VXbZHK/4pmDkQMs
amcCQLx0eqzpnZawxzlS2n/l/SogsoWGuU2g3IH3WmU54F/P6Pn88okLicrinNLFcp5yFZTLhpF9
vtAjsngcVDvP1GhXDA2Yrt+6tFgBIPJlSsPXW9N2Jd6LRs/VmalAGz2j8ejwIA+X13YZoYWTOe8U
9agq6SQw5xABWUVTWMcSuub0gekE2Ui+REK7KmigrZ8QRvFWGrxGR8MDmWW1vTI4ROrBuLiGmIYk
yXMCyqDdvfdj28lJWI6LZKQ8PoDFs3KEz+xK6gzPzvzlyBTOnyo0Xwmurn2a0EdEO53+9ch9RpUs
ewiTFh70zJOjw4uUJp8mQkGg7l7J2O8M5YpqbRfu6FmQm7K1z+dLI4RCiI6yZhF1vXTKg6q0P//U
tY0i1oAInbtpjtp80SE6ZxEf4RY/UXc194yo9RpEdD337EXb4kcmyR61KVKe68zw/9mYmEBh85qf
Z/3Wu/oy9qzlaAMdRMckSAOwuRi2xTo80gQP6/rkiTT2hrsqXkGesNDi9eG3rICtBXiiBuADLRjn
TNUyqvdKaogY9vfhv/Iz0l7Qme2vzAM1AaiQlfemw0LrZrx/m1k2hjl50YqVKFg05Gvqd70XDbe4
0bPxtXMz+alKKtHgtZw4lOPWWrKAC5AzCQk4kyjeAXrSOOxdBNItDgR9aAp2QXNS+oT5Vs4jTIb3
pGPX33/UWJgvmqBtjM8p1zj8YPgSfqLHz2XrJVv1inhXrJ1oKu9aJXj4pbvJAxwef97KCT5b/cjr
HlB4AgNobnJphgq8cgQxaKg2OVUXSIpON80V1I1UxcDLnwGPLdJY/KhnQMLo9ME8W731V7d2Nvt9
3Eh8ivdXgjfvj1DYQ3uhhUeqy6ecUQuzWnJ+kQCEPLR6X51k1doMvRD9uY1lSVShAjDfdonclZKT
3yiV7qsQvak4o0qGM4vj0uH4Ke5WirpCEToc4kTZN4+dyiMoEL4mIJ/0fjoFlV7hdPZJse3TvbO+
l7UrwL5L3zP+/hu0FAVuek1+4WEu6qUgi9lAfTmb66BZ1dFmEsfxAgrdRl+vwbvO34v6kEWLLQF0
7mw0UpMp8tVJ0/NXuDJn7Id3kfbhbZ2mbfU2jS/PbQ2LW/4R1gtj5WfWWWqEM/OZGT7dj1EFd7cX
2YZHgfv5Ygz5BLcutXLXSgrOgWdKC9RelZ3QhL3gZD+Fbh1bvscZ9qPLjGnPUZgWgc3+JDvLiseC
d+1uyoi+h29RC6cUtVmYALqiuD89LmiC3XusR1Jaw/rMfNa+70eJN8dNG+lBkoxhMtn9SBPuKr/k
1+VR/OjQg5vzMTFLNd6+ZiPvuyWiAaHp9j5+v+d0SkBPhGJzGhmf5ykpnIK8fQhxpaOROPq5lHu9
AuXjgEyhTMFiro/3zFWC5ivCgR1gpKOf2NoZyZydtlhcSdySOywwqevPWw3ZhDFtD5eG7YT86nVR
8Y4GgdtfXE4nSD2ow/F1q2jHcWg8w+wJ8myNqHpJfZocsxtQqhsqoHwmy/6v8ep9vxlu3aM5yywf
Y4sI6QzotfNe2hcIx0mTeTwc8SUs5isiU3EOG73DCTzM8kB7Lvlqe2aMTyHGkLm3NZeHSoFHpH/D
r9bL5HvKSjU8NbUfmYynY2+67IKkRgOGWr4N3pVX1PEk1hh+J5V2xQjUOSET6KoJGKTh40niOT2m
QeQdhMPSm2c33LGRM5rsDsolS/pnMbrdqGoa7nAjCzWVWof9gNwEYu9lawKzC3ajss7YGbwiXdFC
QDTqbA452zwFrGtoGO+iX1n64+JtK9PLq5oWJGqnlPzfdDEGmUQTTuXrBygHtp6B7UBOCMOEQP9b
WNXRp2GQbRatMtCFzUTkTkktiHFVhSP5sE36c3uLgpMK+z82gI2GoGE2k7QjiNlsgvS8sfL1lavZ
KU3vYCzJPeWdyre+pcG1RdjyeBiPobilaQy61aIgj77e5ruXzAWykTDSQ5lIINg7lsZoHuNXf/gg
GQkdD3AWwsq/1vnqwUt2RJ7NP1rxUpspKw6NCyE8XIyYQ0vK94dfDdr8Law6W6lIj/SYK2tiQgnN
32HIwP5HUQx36EyrKA2w/I0JJqQ75tqRuFSRZDu/56eb/kZfPKixqmgBTSZrjvZI/wsMASc9Dw2S
1gt/wEHOQjcDeravF2Tjo/kuGC+nh93LYTKkqEzqhjX0sp80W8vCkluc+769XziHLpkKgIOIeDvC
BnSaYlDqCO+h8Yut1GyNDGpbMA4wf/K1nZgihiQ7u4QfL2u0BEsqnKaWLXWzXXWjRYr7Ac3Zxrq0
Sl1b12dLfEi/rmc2cNwm/lJEtVy68dHRFga7bfIEzv1p8wd6LK+AH8kFgVW6h0ppKJU7JcmB2tcA
IEFQtNJFTM6jCRkytRFqoQtTrVzoxW7n0nnhRJkGgv3ROjWhupLkv0TUuKCqAb71RMKnGttCrLPM
XMgG8kVBc6DRFmm3x/uNDmioaMg2jA6YcRAUhzsdM2GDwL6C7UjbOr41L8pm5ECHJKyr/O3kXBKK
NZwn4+SRFBUpSybjoFu2SphlaxK7rCZt7hKgtPEzjCbTUqeUSm9bYQ+xpmijFKOwHZznnARO+aO+
mlTS6VhHDiRPlzgpxkZZFmsvK3+xeitK9fQwBrhOe+kqSk/6nIv9nzXxkRLVIpZaFu1KyiILhJ+1
L9Ut628x47ZJFrW5G5lep8khPzJL2XzHy+UmVBrO5+3h7/4zbdVpeaSYkrudgIIzFjm4+i53dgj1
9/rGc8ELuQKU0To8rFGOZWwvm1FMsY/IQTtgEeZRNCYRhmUxPpvkeYNbzLZRQ63oprPQub9mapk6
rzDIVMo+ZH/cffsvmXtCSvzhVjmf4DIJJRSv/mGzimaJKxif4YzIBVAdk1C9yB7aOQgIq137IcXP
eADxhoJq43fS9ze3gSPCl9xZ0SlshRYKTazXTv/Jvck81MHQDVoJ0qdCmIanObIERREfRaaQY4RK
k1nNIa9EC0Stgoaskp8iSnDHLdNtLv1x4ASz1eR0M0s3lwlXmC4z873eiw7CZSnpEceawmgf68kY
ErxazWOsM99FMTRYqFOFESciYqge28+TcR2rdjDtstdeAMZgDIfWnhzmCh7APFInfxoatuoYWQrk
2wuzNIEFiBCASt8XJ0apnuH4VbHtEJzV6rCGSER4KIGAHifyQ4B3fcy84JWdhktD5fuo9RNLssYm
eSKCBKfd3qtUFIaH2Q9x3GBHALrIFWz1MqAkxCNo003sKsNBZAS6qnhxjB77AnXYjXLGIcCgX0JJ
7nMZ+FSRkn+KoRXoH414lmayQjd1ywYJYSz8q0nn4PWIOXr6j4ksJFq0ss9wa5cQox5T5Zou50lY
F4RJ3sH5Y492bJld3+gsO3PBxOWVjjk/46w5Ob7vx1XvobSYNBY+s7qixjcHBkv+4Kyzw/TSqOY7
q6+HU3kIyJZkqkYk81xHoQ128sV8Ss8X0i0Ofldi2r5td5kC+5e9di6ZcvKhBGKyLTEqezmvCtm8
uTCLE67KonWMdZWZrlwJnwa77JW6VFRtEn1nzkPoj1VqXXr5+AjPzNnYGhLYe/ab2vMq3EOd365c
w8P1O8lE+JRAoPVxUpZmhtTVvGNs929YjTpvK8e5wRohWWonDloCbP9SsM5bEKUIH6SyRNOOYDsu
usnMJ1HgxFy9WQX5M7KSotPRYkiITYQDwJ5iEd6rfsAZWmpAxBjfBwt69hFlk17ifBlWKpSyZuan
+5xlZraFkRo3Wh7Lyey/CfqbxDIV0jW5DXdIG3Y+lxVO63IHwd00iy8qllGMn9AeozYVthLw6pri
PoWHajlhNAwoyKOT4s3waf99Ge4pKWyo1e4k2mfQWY/TzQVjF/PnfFmlPiAp+LOLe97jAzX9vSu5
wGIzSc4KQfi/qtZSFYkBlOhQVaEat/tJdUVf2uSIciWcCBa7/V10ITtPacYqU4UQzGAd7dnEnr0t
m31I7FasbOYK5tnXvffeV587/i4jn6SzFJEQ5z0OfGXONerD5xWXKTK8RqoDoPmOUYXh9QhcVMn+
RurhYbC1GNzvmVRDHvhJlxwaRRTHO5+aJ3xTyosJvBUGZ+ceM9JJGsS6mshomN1IPHdFpoAqkjfV
iS3VfPE0fyfeLg6oKEMW9wmEUKAA+7B6e4MKqWwXZtzFjnygcwWaSTxYiN2ySJIDCpo5lggp+pLL
Xnt5d0UgCWQGTGHp8vkoolu1UHTqhhxenuJBpBghGx67l4JjeWKD8U+Gi2+ib0xz+4R6i6yN4YAc
xK+2LPf+SVAXwzBE2FwTOFjThuYhfPk2OLqJ18RVPH0vPnmzLsPXTyIpmZX5RLpQo8VZTLURwSRQ
GwPePHrTlS259a2svjqWkiDGEe3jwm876cUqGpmHzmJVWFdQTFq6TozpdXTsQ6083TeYTAasvaza
5fAlo3z8QkZXRR4JO8UiwFiiCx+2Xx5Jh5KPZocIV25GQjbuVjkTDQJrE/zRK1rx0ITh/WjMtxO+
2pXjkq1oLzV2+CQNQNSyNJKfakjOSB1oOMzcnks0q0YxVB0Vtn7CyCDp3gutsGQ6P9N1epv7K/tJ
w7OtFre345N4LV9aY6dIgZoVrL5LqUvBDYv2ucsIJM78M8V1sSmMsIclT2HdMax7QZvnfyrGsfKm
Wj6Iu7o5s2er5ne1bHVQQ4jfrmml4F3tvzNwX7TnOCRsI7K1BH2pID0lIkF/stMLqfmVphouGaYz
COVtGHDzK8/3q5tfd7tvfQNpiZQrt71tUTq3qW5P78RXohkF/NrCcQu0hcHJUl3iUBd4lmKIuMQJ
vXUu4sppG5lj4JXfCePku+/A1pBeAmjhCOtEj9foAtoZuw+k5VNTdhkep9zrqCLEu9VZWnEhKu39
wEGsEHERqERqvaiHBl4olXOhGZ97KiCin/Uqt+uWaZWvxRL6XuVX4iohiIRssS56+GACWeMIVd7/
x8flh6w3HNPmx1iTCEmhPt/f7UIybg2NEYteimdaiImE1qSdNH4gkU4mEfvq7+bVsPDMvV97J/d4
LD4vikmsujmkl/Sv+NCRIybcnoO6IFqZg+xXASbou1TB8A3ern9qXPQFS9FA7rcIE7NP8CQIjXG1
IILYTOUVakywvll/WcU6tf5lJXzlHTvdG42slMG3OqQJAHCvibG/S80gndV+HGv+jKnWsyOolxzj
WikaK9qldkPNrc8c8ceGKZQBRlXbzK8dbrU3P3v9UZCFKZCc2io81oZqgJIuK2jORhQXIgwwMQcX
qM0kBMgkRIS40AE3IWVZD5Lyjx0c7DNJuFpCieIx3K7x1wuU8Ki9oLdSuux5iVLNG++iI2eYprxa
oZ46yhmwFr17Jj1faztghreKdsWZEKVTSGaEZYcRonvLxz73X8GwIn6eIyFz8cVnplbpyEivCSg7
X4FESVO+V0p+BCmwnml6wZ94tTbBKdKw6bNwMCa91OhVGLrFDg1weNqxClh9TU57jWJDH/xnPZ4A
3b81UA42IShmT+sCBrW/i7MqwEdfJ3BMcN1noyN5EjqxJzjq827GrgZDMNMy4d88PIXf91yleGrA
7gFpXVNzS0MEsjPAo75CdfLHje+/hNy50jRS5dNnZVHr2kihwEzd8JberthG1/qsD+4y0dgCWgHL
le9x+lEt4r+rf2JvxfgpPrjCbsj25peP0C3TcxSdstMPqMhSSmOR9TpWVrIfRbMmD2BxHzpKXlaH
KYhX+AAfs91clRFeeFs0X/9rPRyengIGkJHOA8GP8SLKcCwNKj9WqUudm4kV0+BJX5kXsZ8z0Dp5
ucvcCDN9xamuU2ti45ZmCzN79VUslcDDN9sLx7USQrHGBJbz0qKh2JSNXoLG3jxMldx4ZWFkqS3+
1ys5jXbaot1nwp24kLKaT16G42D/4J5Rq3UL//1AUUlU1K1xzbxDfKMRqjf3VrR2b97vU3vekGUL
RgooOIvSFxjdzs8m4fufJSyyA+k85IY9DbIu/UFDI3QRhx/V25kA0xctsf6NQdxXYvctfT0u4C5H
1z3FnoFcwhqe3n5iZ3d2VHsmmgWlzZ3nGFnz52CF3abUXlEemCSOuj25kLLfOJLxT+83SGsmbaYn
1F/1s+mWJ2J2T2RyhroSezlk+5kgLppfSr93a85qsYrTr6dxgLtpESNBP2huvAXb2WjA1vsAXyPu
Sc9a4mPUgIhyHOZ3JlI8lLecY79cUNlcyw7Zp20iNFNqjOJB+VhBS1uQQFfyGszr3u2hy6pKNosh
z5jRb0vW19kuI2PJbAaD85jRjn3CJmNdGkahS1wwHW46BzBH11pHZHO7KMZ7lb9el+rrHLI1xBB2
bG6D3Ivgb834FkCtGMTR2mvCOEWX566gJ6KLUJpD387AYZvNn/6yL1wnuPgPArNAxLLI0WJdqm7Q
Obsw31zaNMRQ+hZIh3ZxIzA8pdEMXQ1JYQM+b2ZBRRt5/D68MfNiCfHPWYiOjfdUXZsLr5Q0/mMs
DuDhyzPTKSdjNMP4x6F6/iZlgqqUEGqbwGGbAl6XFQIncdGlZJhXAd4Ddui5kqrwV59A3DZgbIDy
9jAzhOV+S1cmwFkZuVpynYuncZEe7teCj4WRzgXk3IVMHyVBJ5b5D1nlOWHysEpOlX1bOItL6M45
4fln3Aehx500J9H+BGq3487JO5d9z1JYCx9Z/QATZeAh0qinSyUA68gN83Mu/wBRm6gmELni6eYq
im56ba044qKajR7K3O/9lwzaHj3rzUSw7owxgU/FyoqtZFNXl9Q6S9f2/ogIH/v33/dExKyrN5rv
mvVJVrBwYRGeiaL0cmYtfwKo/RQ+8TdSKWfuAsx3dI5wxr6nHB0UZFSoII/MBqxHGMk1C4pEq/ZY
h1YZoY6bYQ80lZPJCDqOScmdgIgqtrEstaMHF+To4piZP1lTSXBVaKnFCCc93Uy8N/76dmXYa3ZH
2nIQaPbiuu+ricY6xI09zfLdlMSbly7GyUEv8vLZsRSm99YphNjLF/IGMuqfCXJ0BlsqLUKdKiMd
4dYTSrR1DoGHeau+CEnQ0WqYDofN8pHto4kQvOi05Q18UapVG9zsFsOlUHXGoNkivu4ijJcrXyos
e+s4031F6ZViyMe4k0V4kd+mm8FhJGzIzPNqw0bQqGdhOvm/XVk4Qw8CrPPM5aa2F9I2wMVj+Bzy
pYRTYD8LflwFc9f6q+m0LsrGGU3+Ul4PI9df+RC/IdUkttIbTE3RpustFbdRErpEw8K6HUCynfgU
BrsCowysAHMJEtVD5Hz8DQ5pZoe/QsYBG8pY86zQr/LrRzmmaD3uvrV3H1Mn1+vLcCUJqvTZ0GPR
Q7EcyMzlzTyjEmUFhIAf6L/ePIBWWaaiezerNAfI9Q+skJ/TmCOouxdOnnm01FQl7dCgV06ziUws
Lb0oIwEuwYw602i8htGN+yKxQy1g24lLIKK/zp1s/sosMRcWgptLx4PadcjB+fEAl7m3b1r+JWMI
PDFnniJy8RqFXI1i4oNDd+gIdYQbGV4NdzaZa9UjXMvDOs84t9VlSWKZTb00Pl/npkK3+PuAoAym
uH8qmmDuhsQloqzPERTykWPBKMT0ck1Q4AwP6CYGRCvUYwRLEBBEAvxhxC2c7FyRgcpW2OIaRAeU
aG2LEAtfTjSm653mza8Fk2KBa3RwW7M8MypJ6+wWYRFGGLIYcf2L/G8TMNqjUBC1d+IeIzaimhs1
ZW2DJMaEgABkmwpnrSH/qtcR/rLtlgHvd8/H4eIg9fwVYVfq2QtzTyYtZf5dzaD3VBsllZGuNWGM
DOnT1caAO3gI8IV3yHByIRTuht8oSZsdxSj2l30tuu2TyAKxv7qp1oijGN9haDILxeL966eDmcxm
+wUKCPKeXinscXXk2vURbnHJJjaUqxd2JjhWCkNnhxxUpn/ARAlPDTW35oKJnstKahR2vtXvyHLT
4QwWsLYizTJ4EHgcAIok8nZQH7jicELHzfulvDT0JIi1I0EBC9lJuEScqaug2VNt2Puh/8nt9XI1
q4OlEy8TdquWcrdLgwkjUN3X8MrHSjY1cB+8ngLGvm0bqUR2+E86px+KJtyKCfi47VuK8cneCGRJ
zYPPxichxtAOQOwRueLhBek+2EE9yYrNZ0SOUw83f0Gt18+ZD/bq9ysJK0v/T0SorXP1z6g49O/v
zWwPpRJtvsIh0tEe919Vqlaif2klc5zLrLIYyM6Ln3lQVcR+kqRPXiAUizx0RZfQ4QNYhfATKeN7
WZMNvfrmv1h1wB5HBiLL4xV8tvcWzAxgWWkn0U+yW/FIx9ix5n+fom/m9Zxitd2N8a+2pmamCFF/
cOxNVnlf6jstyPL93EHRrE3icVaaMrBvuhB2LheP9DkLEgYRckqqFnWSGsW5pUr8fkxL/FDIa5oG
XjFPF1fKqicxXXtrmnTbsNybHXCKIdn9BAs2ncHPB7LQgZiV658YC14kX4JkXveOjtHB6QVKnOvC
SbsuBdMxIdgW8J1BrEBxQA1dB5cLp4xfzR8E1DHxQ9P5Bc05N4T7huJj+NjnyfStxqdQjvu7g03r
H17OkI4mFFzFAIXiyy/3RLuVCzSCxy7BBUnWSEbZdO76hsmreKncK1YZfjdSpAoIHRwEwNSGwgKP
lYVOXb4Q6EZxTjxiimve65yJQiE+6pXnTvjLGGtoXAQppfFQP6SyW0UKrYhcciDBeIDmr9b4dNAT
4OLyZmAIqEgvZf+cwsE+EDCTqwvmb6sDhAHtGrkZYxG0PcwaD0v+YLkzG2lBVBTawnwOzadW5Jps
othLi2xcph26nNT6kROg39qMj5t1ecpdVHhheOKuMfjYaCBwl/nCgxW8/kncSHyY0YWnSNzkIbzq
sYpdJIKFBIDDBxxd2ueJLwzwueQCGkcJF6nFAoyDd5dJ1p4mnqFmWfhXcu94EElPT2vFXZXS1tmv
DQsLPtYjTjs3I9Ft8zNFR8DLe4IJMD+tvxZNPuAo13JahK4Vgo+CJi8l9JbE+IG0NhWCW3M2rIWL
8R13MW2/Qs4vV4wQQ36o87uFXqPnDuN/+ljjHqZHKpAbRtMkx5xDqYB6fv806WvwM+ZluH1JHz3u
QqDYrr2Zz31CNWqdYhFv+bwAT0wcuoeC8nfPyr/bXIVgwXSACmtKxF8mxJgXvqR4hiXF9KjpU4lf
jixX3ypHKLctbl44Yr56kEyNtn2I+6bmbVUlZ9omQpicfxoE2/D3Y1qJG9TzWSf+pnUjvebHF7/J
1AZ4qLlsqCzeXGLlhGCHLxhYws3IoS+w29ue+lsBgh0G0urau4HbaKHdfj0p6iVhVOLDgQs8TCXA
VdRaxyIuNY2SFYLEMPFOKsnX8T1u2JRUYzt9hg9SOV6NrX4GEdrGh72wgQIRRmFepuv7AOf3jls4
8j6a+HXwNwwJvGHnoKv0ux32pWdgXDK8QW1Mi3gAyclgMvj4g1K5dVwkC7DqvFL6V/Er427EAlCT
5Iha0QF+t0UL8H9zBzt0Sf0MlrCHHsM+bi8LcEoa4eiYmdtlhZ2PvBNqOoOvjDASDAQEXNwkq/zR
gpkVPWvQBopka9C7rb2w6hmiHcm8UnyjBW4Cezb4y0JQGLCMDR3a1noqJDTsZt8Dx3HhZtOXibnH
wuUAgc7NYmp5NDwfXMX8WazvT11L4K3IEEMD2MhE3VuAl+gzMLziPI5JcZfKXwFv66VdarHipfWT
W9usttwhi4dnZJTlePTh823aYHaXDD/eAG0xI4b+LP9BuWip24xJZeW368aM3Au/v3nkoQjaDMHE
VSWogJUkNnghLQu29r3NtjFPzSJpgtvX/CGoz+x6kBexifgmuJn2dJxZXR6dyMdCr28u6BxNVVU/
NzdONo6rBZ2PFKt44UuqnTmpeHekmHx80gUHHf4GA9Pm410hAeyn6LDyAqaGZdPnKXffKllstApR
Y0SqkJQ9WmrffvMJbnvEy6Cx/g8X513ATzd94RIOscAp/HibuUIOMaS9uwFG4J4Ihqsndixztaw9
Xok2XEyO58VzVKo57/NGwHm9HBBAYifIlTp2wNVrLTMd5XYVAujIwtwSURMxH33jknOXJdvpOzEP
KfjR/wWxrzI1pBGWhkDPu1soACxVHEd+wX9GN3z44d1ETTusNakPyyHJbpxrKZyHVvA1+/walGLr
UmxLZCUsBpjUIyFjTUQtpev8029KQ4Tbnd4c1NmvhQUzGAjRPa/rMqa3GTeub53TkFuwiCOIenHw
VFuYrMdCZ9Xn+V1nHtiYU1m+HfbLCft9XBCLWjIRfY2EVQiHVgtyptCpDzzEbxc5NGJbk7lUGesu
79xDlJH1HeuT6CjlgwcWGbQp6Sehro1LsIYkObGrVOrLTQRwKztCsKGWJxo3y53uKkjMXF5tTFEF
hxZEOs3fDecDCT23KOLONG3vw16f8Rqx/4fjDJow8ayzuA0u22mOOt4Z6GkA4ZroPKh2/cEfSBKd
CKILUbH99Rh6Gc8gwnQwdAQyEmPHuuZOOz/L843Tb6sb5MFXwRo61Zrxzwmq8h5m40/iVB/aN8Jo
VU20eBYgHH0N7DcHIQrreIyUweYeNmRSkFU+byzoHn684RwwDfKqCTVkrtFq5IydkULL6AYEKrMB
oo1PTcFFRvPyHNQcLmSUWrekbxZ7Q1PfabsaWoEpeGvrIghSSr5mMOWoyJpp4R5132QK8sZ8qQsy
3vXs1GX3Ja3JuPh+Anoh1s5FsuH7doYN0bBb4vbvh2Z9sRM5Go6IvNgxEEq+W/wxx5mdjdiCamXi
6zNkAeFL6m6zysB1G9FhpoSHtXiDnAMkFC19svkL3MLrdtfm9cwUbSiReiQP+w+Yuz96QANAS8xy
P9JlPwa8xDuMsqoUdPFN/6eLNOEvMs9zM8s4nJ1lo1oInDc89/vBNjN59/qXyVdCt0F967e965Gt
trAwMpPrw3J3b1nkyHONCQrPvrfhBu/FYGmZ0X7od1JnvzdN7/FzobEYHjav/VDmNrAax7eXOlpf
1Epo6IQ9lyBx5l79wNcOKL91N7VY7JgosMP2IZrsh2yzasdf/xVF3a+NrH34jxE+USR6/lobVwoj
FtpcEHRHjqhckXRzOQw6n41Icovkehgc5F0m/0lsuQ5XVo55HqyX23uQdX8a+Vs2Y0VSs6/4DjCo
41iJonLn6v3UPbxvij+ItsW4Zwm4j/U=
`protect end_protected
