-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
boJxu6TE9fXYuPf5ajELC0cDcRPlUo0hSm6fLyyBB1znvGIPMAF72ikihgcvXV/y8Rh0DNRVUUQI
u13dJQGlpYdVdeo4Ln2JEv6BjNC8omFAR19koMt4gFDwGGkjh9xWg6svJvw3I2tGh3M51opn+D2q
OKo7URN5CTbnEAK9PjHsvVjBz73UQ5NHIJMyMtTsxFptsd8VGghcirq9YlLXTnHNgIaFTSjLc0EW
mXgauku8L8SrXlPn6BajStty7Z4/4dpWjPW0BuJlNIiWkYy7Xf6s4mxcqbVRA9HY0AEzbXhJ6pqJ
SflpltzlHWlbHgSmVVGOm1qr8S6JbwOXltx5NA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 1072)
`protect data_block
t0cFlEKZAS1CbTwDqCEEmsK/wBnpNunKhbxiIluYboT8aNlZ60R4Bv3v51joD7CF66EEJTyV09Uy
lCP8+Xcnx9zYIzSZOjELTQUGdoUnRzSh092S2swvawriLjmcvg5/GMYuvrUj53pPLxs8t88TZwaE
JVch5m/AhRn038wyR5GFzk1hY/sk8ANgEpohfTHRKvotO2mxeURnhGZWXsd41v/O1kEt1dqIIdet
wMwBZYb5aUXKO/e+AvqvSpWoH5xp6Bbe9XK+TJQLUbgeOtqhm8rszXIvJZrcOzQpr/Is3vJdcr6D
e1sa0a5vbZ9IEgqeKTYB0PhOPu/dn2Q1AtCyA6YaxRsTHPVlidkHZyklLwIy3OLuEO9Ue3wQu7Ax
LR7ffvkGNtCwikwdVwwYjEPQ8skz5TljQvXt7j3rX2BV5qSDu+0Csea0PYrvWmLdcea5mkoEtt0J
GfLYUJ+SqEQ8YVIETIW2qqoLa7Go4+fspf/O9/WSJkGPCc6ags6206uAURjVM28W3AM6tZZTfK7D
ut7X/H4wizz9bzkWalGbVUpxYXLDfx82VJjuo6BRUPUUh6L8HYAkJttx5/6+PGZmb6U9Tl4BdI21
Ar9cgxcfbvFvLgGL9L5URez0htJh8M8wUjr1iQaZgfJAFUIv6ZnU9lL7T2pxrjwCV9kzuG82q8Bu
rswihEsI1Uy5AXtB8aJkd7UZ8nRQAuKqY3EWJ01cmytv9WZ5Udx9MLEXVlyO3MGVxf+1lPh4lGZL
e7LdWZDVhItQUkBUzdMsxtSKbo4uM+8A0d0YpRWR+uAZpKxNr4ieyXgcEjP7uSoFGffE5co9yd/B
ZZU7Dug5AxFvqCxk8IFiWLxUSAPxWAFV27I/qbH+aTx3EJdvhDoZX7Ra6Qrx0VhNNgKA7bpKMnj+
NGBDxoOF3T8DfVhEBX/PWFNfi9ad5WSOeL9jXb0ACYmyNmQgHUC3manqjtcTPpxGDwN5GQ6gwsLF
nzu1s3rCJVxss7J+Ke2LBa/n0dlgRGP05+FjaMShYZLddiGv/7lhHUN2myDrrXzQr2y+SqAi4sWR
fdd+WAezvKovomNyR5zLLKgWTJBoGTJDygv/0NPNhaPFy8Unq+GcnTmy9Qe5/cnfsvnMAWyq4FzX
k0p/be+qNTwk56dPA8ifQxWlPJb6XDfmUZAT6YkLpzb2fL2m/sJFiKChWufCtlG9za0rpiN44/Ij
CaxCZ0MdiFzcTL8D7lD8qysmumAtrlXZ62Isc0ziYYmEHyOj+Ai5SRKx2rzz+mEkIsVSXFpM4GXt
qFqRH2/5H0Mji2XDfGxQarKDVqtGDrh3AS+SqEFFEvihr0H6sioWV4fRdPf+Xx3PI93CkJVyZCyn
ax4kLBOwpDCdEfrk6a88ogrWfMQvQq1R45ZT0zVa7dOSvr9MndcbfZkNdkSS0Q==
`protect end_protected
