-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
VoUbXt9czBS/hp/Hu9WSyByRDYL7yzaya/XDPVEcj3JOKH63oTgSpgc91XFrrVwel8kfaKvirpxc
K22s4eT8BM05/9HzsxkGNTW1FGslvaTRvfMWjylV+EapwUoaw4Jz1HtN3TP1vKYFCk75Gva9bvV+
6QtFLw46ICT7jInJDalmdX7Ck+5P5zpHIbbW5OtNj8jLavp31IQwzJ4jatUZ6uBmYlo09DB6f0Wo
w1uOLnaxkLvjzFSdfQz061hNEeQVQocn8CskXh/4r2HRzrNvuvg9LyFeRtZXZOJI9aNU2NxWasbL
MiUtnCM2+U41xGM5RLADkXADD/KtEtYBcBhiEw==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 28512)
`protect data_block
nBMNtQhpeq7bXOSg80GB1JNSdWOf1dzJ9WQKYGLhnGTopt1CwrLVGJMWYsi8MmNWVEuElqv/0lnL
gRYb+0XE4q7pnVdu0qxQKM7tUT1U0ObvIezCKM7wWnyMhu51LBFouyiBx1JjU2RNTy5GeSff0kI1
TaEhpYXFQaxgV8SH7X7L3++4dUPESygPSD76jvbL002H4DeFNjtsspR3q99q8Q9xoKHw7XlfLDYP
WQBP8S8T0ddhajYaIEcSAC38WNkFQ6nCa1EcwgLpbRo3L2qDWWH8N57+EvpyY8NngKyxEJbsILEY
9MPzgb/F224qKbv17Z+ArYke5c2VYMUaisvnr2UTaziVz0CcYNf37nlCmJafXXK8b/pCMYqCcXpU
0NgBgH8mYoxy06RWut0aBEpoB/FTGpNAzx3+hbkW3tODHQd/LNpRZrqo7DoQPlsDndmSDgFV9Pbi
qPXxFiow3kbMVn2wZpU9+9I1thIGrDTwx2q996/SlOcG8TlQ0Z+ap1CWp5I1Ukz3FJ3OJsy/Ja4l
mS+nmnVGAle7U818zIs0dL5+5JOr03AvKTpugQxCY8ecmQQGhhTUFiFib79ts338Fsd+8W1uyB31
wYtEMd0Tv/acY3aocUg2LvKPpWq5jAAd3q3lx2QbuvYnpV7tzH8a63Ia++SOWO8mc/EW4Ulq49h6
u2wKRAPW4qqccDk2fI+aEtmUrMo5ft+4Hu9gOO0H2CkNYAyPZwRQGwwNbK1SoIACToqeEP1QmxxH
j3cAlxlzFsSCniAr1Ycl+7UE5bGZihG2x0ETdeF4FcGQR1ZIBnGh+DFfYSp1EKq8X1I2cjJP5XUT
S/W8H3ZcXkZd8rGLnu4ickoZwqGNbvptUDEP6DYXtcmVOWM55qAdbxl+DRml+srMwLxjzQ/uiUCC
SZuCqgBSwNLexKPcCtS3g5mhNvyRFYflYkjKVau5G1aJo5cSDfngSejpiSNm2cxml8c8CWYBDREK
buhMYpUxUpVHrd6DuPg51wPyH9JtcOuowwP+2oB/oS2Vil29WlC+PaOUYkaxPvwoFYsjPAJLXOUv
2RDEPS3NQTbaRp3o2bFN2Cig7S4MPd3MncglrZKi8Wi1r/xdUnLnH1cLcsBz6qamxC2ZHCa+6RnG
w4msQY0xDVjuvkDuy9NvmNmRdD8Xc62juKSyKC4zJffakeSPiRnEQ1Vu4r9KulzwV1KX9JVNzGQ+
y21c/P4BfK+JAZvddRy8I73mbMKoQ+t10fGo1pBnBlon5S3dy2t6NNlhXv26ZAyPbqlrpvbJ7qS1
mVoT1kx5mBhPWOWymiDbLDsgat9I+yIE4NG6aoc4Yo4QSS5UTSxY4SOTkhvTq3FHQvqmFd86Jyn2
lE4mNHA/z/fAsFJCWfC5jiM2wrW2caTfRPLlkQEcQjAIUzsp3msdH/F19AphNDdFNF6ZFsF0ZW6S
HCNBSeRf4Cr1po1+gD2vtG3KA57k1DOJ2jkv31sW5r13Ub9tTedxZYwxXQfD9IAPKCHVUOqiOeLF
oji6t3ds0a4V67PrdT+BF/CfJo3i1d0viOcvSxzFEf/rLzjv5W3S7+ZD65whlYiWtA2yh0rFqvio
vlThEMBHFRY9N6PRUU1vzC7wwrXgspc5UoLr99CrgZtmH4s7Kbt/lboatVuzBeRVM6SOMw1jfK2B
Pn58uoJQwiVJy0BgbM37eM2vlPEmD5rb6RC2Euo4tzFvDa1pM0P8H1qqP2Tw0LyHdZT5tXVpr6w/
uwf3IdGfKSqETdyKKOjRMewSPUrHmTfNibfZTw14N/5xRS+0gAcWTJnTCn6MToYDkf80uOIYy0/c
Aa5QlCjyVS4Yv6ZzxtydClks/8c+/ZYFqoz8NVYZszdxNSUzNUh/wtfTLNs6fufE3YF1V/svK4CB
YkcwigcrkU/fpdjenNxiNKAzOxqcZOxcca2xAxOfBrLMPHNjYAVMSIUrqCGT1pj9dnoiUkVup7i2
WwqRxmU5qsc2kgAsiKqfJS/dv6WYIHB8zCOfQtOQHdGad3EylEkgaPMFo6rEaEr/SqvRJFKGGVsN
UBZ93ny0y+JZeXnKEzSdOFFsaMUKOL7UlJo6RiPHVIuGw5Los3sIFfQqSuHNugVyVK7VqvRVGuxi
0EtP5ZOo965nQ2fVkaFbE39tu/FYs/boSHAl/uPn93lUjPXsgWK5uNBl5WncD0D1dCmVOfng7I5a
1NXCNlQZOQJ2G1xabunS98kXcPGzHqe6LexhBCbU4vpg68/SyEVDrItiSM4B9FJBZYcrw3km6FPZ
qajvKzWlGaiFwWRasUVNw9X37QCUJ7/bzd/vTsXj/8hi16joLjxex/UpzGv9BTWwQmVWeCdWIuo3
trN/yqbFZq0OTZ22KPe0i9OZr+qEhlSUeHvRuxfE78zLKdcXULpT2cEMs8YjbAA/buqdPBaJI0EF
a73Vv+L8guLKF3G68TnoB1Zgb8lwYNKrdj2HAWAe6vj+kLBjMdCQLp1EL85iAXWm+J4+lrV6oudI
D1fGMcnqXbXJVc5o6kosOHrF1UZ5kd8AbVDW0ckuBPK/yosTOcUmrox5O61qYec+5H+BXm0GnsJg
kQPioTkeQcLbTbeUpT7jeFhSWODQJbRe4A4h6qov7Gw1jzsN9MSuHfJCMlDcrqd+4krTIVPqfnmM
UFvdCpO5LwCbLHxjA3x5N9ayCy2QVZOoS8sZbGZPVPMxo15Ub6CjWWmNss52ZHKXRQl3yPww9hDr
YPWrCf6b8YuZQ6/POHCo+NsA14CLdMv/yLbb6+cWm1UDMHlSlO+EvF142hjdhLiCiekqEL8pqbVI
+FF5lnjDJ6+aR9R2ImmDL+XrViW6WYBUjEPuIasAotXXwHQMcE+bfX64+O/gN/pLq0I96HC91Bdw
6VoajoG+hd0bMqFzXbKVH8ZMwdLbFH+h3n9bzyKinpj22pSCHA1GYlzHgb+sMvNKRoiWg5zVbcIC
qBZIoDU7NLg8OgZ8Hdg0X592xpdoAQ+xzmAETLf3tcAWq3fA4pbbhrrk66c68JobqC/ljNe75PEr
w2y8zoXoHgtf+C7FoB2HwIYmhm5EskjMpuHAEysa9ebY2taJqfHK4IUc+kzVgFnFLeAyUQ7nm3M8
9O1Bd11LGR1D5oOntRA+PhcoI8dXR9Ce/J9m4xFNia1WOQliotds7DxGJUMrcsiw+mW9+tFt1Alp
CVwLEn4QMJ0n6sX2x3MVnHdkWzVhrc5oq3d8I51fDL9D9YQjwInsrlb6onAS/+LBtT7T78fvy1tg
f1q/R8YXh7im4nsPjbePAmqxyinv0g7DHzvRA0xWTYBgo3nyqyYrZZE4gePU4GDC7QS71mFX6Nec
7q5VKdjICX9cH6QEv1+S+s8cou5BbqOH57as+oZpTRT5zozay3GisDyhWw6Uf1Iyy396Q3tbiUnS
kte67HBTV38ikrvb1S8doBymojbbdednQSJx/Q9N7N6MnZbusjgjZAljXKmnyBE02Hq9+Um5+w3Q
MCOJz+7ketkTi/z0E3ygvWcVS44UzmhsYfbt6SN7OxJOPYhlPYEvyoFBpE3qznMgKrs/c2pfmVnM
eHj8nlg1vca+qoFE8KVMwO5XB4MRZaGUDWYxu9Rg/0EWzfbqT6Zr6eivLHRqL+4uwjcCEddpw+vJ
zwA1tL5stcER4Tp3z8pHlFApWsMUL2LPlxF5EA9rGJ62cTk1cwDs8c2ChgqekpquVeNS7gCDXAW6
L8FgLZtC0ASLj/KEH0lgRMSjwOqeDuHXotfhuUngqlohOLNXeX3AvAeWVDmAvsvzEM0V2o/lLosv
AgZzTY45RvJMQjBekwHTsYLsbLPm1cQScWMzjAXIecrJhKSMP0djjz5aQSz1ygakQ1kifnvjyVhq
JMcbd+fUyWklgIUtdA61B42ELK5MueOoB269LTxiy/3JFxInzAgIISADO3W2bu0Y44ZkUV/2MQ8X
W6ycymQNIlM4r8c30Y5VY5htjWRaEIA6gOP5e5GHIFvyySZv0VxHyser1S2s4JhzFQxjZzCh1A7O
S7FJDcI0esgwz7vX3h3zDGwO3ow8CwBUbbhpVBuiQD9r/7gM0NRWK67Iw0lJGPuE+e8GW+toN8dc
mdM1GSuGa41na4Izjn/kmuzJdEiG9KBhPsPn2hhPkxZ3q75wyn9rCCOkyStQ1w/6NfVvPcOB2Cro
6lC5eGc3+qy02qq+zJ23pFfV2boz2r+YK7mtZCxvjJPj8Fyuy+WnHax/P5IJBPqnYTMUfzt6FB85
v5eYq95Rn/FAiyDRyAtH8EyEAgW9bSVKZoWDrtH/kIhg0G5AV/RkM4LQywcpvWaxxf5DGp717ekL
jQA9SzJgGH5DXeDDaGKmg14FvxPmnJZbBDgw1p49bBuaROiBxqM+VT9yG5SAoShSG8g5Oav4LgZV
no14bEc/axDiF8aLmqM4FqJQPwAE8zFPvStl074aluzdLYoAWZlO9Yfa41n+iaXI0FUh9oQJbno+
VfTGDK9h6XY0klLxE0NHr77jqFmJhNoecGR8oTOeWPkH0oj5aiJRQwk3PkoigMKhHausqnNQHXUs
fHZ+sW8p60aYssY/SedUHCWmqF/gIexFV/d9EcRBlYVYpX2C4gC6BSbSVDBvFyNR4gcYeEjhWFDi
bWAxOu3WQ2UpJoqZjD4F458YnTVq8CwqhyT6ahJzs8oWgjVjAdPXN8FAbqyt/z/OZopXyc/XyNw7
MXdx5BArJMsMcP38aaXADkJVi8IQVvcalpugZzgaUGQZUUqJAEbzZAMbmKggd77wcNK79n3XYlZo
PaZ/NwzHuWK98len3//4riSNjRauCe4LlWuHD/iFdle2uugqh38Hq0FdaYSKNCS9Mpgw7yL0qHPe
uGNG2nfEZS+t0iTQm0wceorMGDpvntjTQ1VHaL4NahjuoT5KXYyL2LHBFG1EcbcCOM//Mhrj2yPY
gMmdjaq+XmzopvomLTLEIm6E7Fitwxo7bAUdNBHlg+L6V08YoHYUIq4lObLWgK7X1XfoNORUCVTf
qpaKtfok8tUNTvVy+h907L7LqvArQb9tk/PD5cV3Tg6CAlPrQgb9W0Knv56LeAmoi7EVq0tQ+zTq
0sSseKH79V5wogSfVZfYbBtvbOFP2SLNNfi4FlQl+MDl/pYERD8kagxogP7MaOoGa4njaTYv0OES
fcG2pflnnqu/0Fgl5gwXGUcIJ+CO2gYlsDdyJtnVfeADAUswPKdxICK+IfPPPtlRQMUpMU1oy65w
J4CDhkFCmgUNLlO7sz5eGQ1vM07OVTkBBLh5CvkgXy/B/lCCuTmNeelA2AjTohx1kqCxAeMtcin/
ojBWCFqFIdZ5K+Dp2ojsba/3zDtBGJrzyBIqkaEWk6OnsxpQJIjOb3N6OCr5+KKoDTnTYudE1xsw
4g895elCNMuYzjvXIFDiPXPfZxQeeS4J3cwhHmTuyLga/BfCL9Fs9Q5X2pXE+lQ+eRcplY65pDvi
/ms9R2wwOq+mlP9mEd9VsU6KUAV5jziS0nTfB2CApFsizeNReBmPaJmzhgVU9pR539jipgNLoRFU
2FPDnEhq5G3TTIh+JBy0Re9KEVhlwpMFZCCoI2V4lplCWmpDxN3sdvB8pw6zYCdlx+iwzr7i/iIN
Ghm5WyVN+lv2WvO22fRAawncPR2XzZvg8v+k0++Fe80XV52Wsm1UetXb1lEtUmCNHV4iOIH9B2so
B4qzGgz7dfWtY0g6WmzdleQ8j5qPslpgI7niRPMun0IkrEyC/nKOvcO0nmSbHCf0LWACTfDvLepk
WYGWFdZbKmjYZojVhtoO3FKxZlnFhOBPG/3bzv5r/LPMzxVa0X2+galqRoBmi4ngwgBTLLix5W6p
qErKBiJa8ESyex6GxTVo7kZZNRMo3sXCOwBTMijeH+7r6KBBFhroYqodGGbmUo7jHYuX+I4RHfnP
rfiDkms/OKVmLLxbDy7J0jc/DpjT8XXeRntAOPaLclfb/ro/NXLs3M+OklH7vuYzZZUTr9JxvgR9
TzEzmLzIn5ZmYph0fEvfvPT6zDM9iJpvRgAXjxySwbGs++ln/4L+0RNZSw9YKSKDd68PsK31lYzW
vfx9i4WI/Bmn5cLlaEBkS24opV+jVgfpWCwRXx/uXnYj388Xw3ociUC9iN5zJer00ZZEIR+uyQuL
6dMpWoD6X6jcCH6/yxSLjigyhVXoJX3ZD0MQ73W/9dmCQZaPqMEY3RmkpnQI+OM1sE2fPnKYFobp
xi3z4joBSBU3D5sB62x1U30FIzZb0wlKVssw59XIHTVWDWEgdUYUIOiAtMrvEId43aD2pKTmPAgA
1r4bFLvPjpyQgQsl2hWYGNL2vFsR0rvBN+rQw4UOLosNMhz6WUDtJD11vz7PjVHyc0oU7Py8Lv4P
ZTE0dV/1HAjzvBUWCGWEXQT8cR1f92gSCxcoTBqwhgzHmfSxPkp5Kivnz/Wx/AIMsrGzr5a01zh1
rqcay/QIylKEvTFPYusoHhrObZ6fhKaTebYPRf8qRXng1A6KxvJ7/ImiaGAy0vM/FsWBS9rgVupc
VivO4tH3dikrppvxq5rLg73BS7CAYPm7G6PUk5fe05aDJUHK7E4vnXj61NL+caWTXO55KY32dC7J
mqvvXdJdCIeTmFcmU2QUw7M0rWGCJAg17rF33VBJF5lYz0yjWBGuOY0pEZgU3otLBcdZmm2vjDZ0
AEQyQ7xns8Oa3A7XuU+0uNBjEI2lCv+HFF5E1n2zBOrtFmYEfHTz/ehkLaUZ8Mjq065hXCb8pl3t
wyCCCZM8B/D994xo9Qy579LU2zRO4DbzSm2wRjeABw9yIUcjk4L72KiPOPLB+ZbVNQSVnNaMttM8
gNkicYTFIb7ITBeessPZV5YpBLWOymsk/GMEtH8xniQdxsjcxY/1LcdMiULgj3eZZ8Gl38Yvk9eu
q1MENZIJaogmH4CDZeNSYUsCC7t9+4IVQ+bRJbysdHTiusdXlvvqJOZZo9E/po67+mpExEebslFJ
nbSj/IxYm4I/hitQwiaHPeBo7Z3VzNL2SLIJehvfEWvPm825iFofkNNjYECvBJUZzDD/wiY5TKf4
BJIS5YPZp+mwNZ/hH+OW6EPqjJu8tf/TR+CFGG8jvQ4MDBYCcnYJZGeKpiAbQA49CmmPJ1qepNmq
ARUeRD+sj7RH6+yATjXAj19cX5EDRVZmfbt4UyMXZrAYcImAIDDnp9dSiLLspbE2axavNs9zCd7g
FyQ9T/lZ6dXP8mTym/TtQFefQCOu7nwqxQ65VJeJWekbNLt8sQBF5RKfDrxtKZ27zO7TIinBpCTe
zQEXJWbj+08R+Y1iiqScO1dzaLNwySAX4FJLGZSnOhp+8R4zg3y6PB8fzVIQFZbiwrm4oXJnlG+Z
fypdOIkqLANfln8uZ7tKAoqpCt3MI2lGnPFfmaovyd1e3Kqn35g8NTBd24x3ZnQk+4Omf78a3WEF
OqLRpJ17PE0rrQFTDg3oQsTnAeeRbR4yJ1lfMINfKptF7nqV5Bdq9aKdVoa7Wj68E1QZvdzjSqQ+
2KUrB9LNjiL17o4bdolr6VreZt6NrCE7U1q9cd8B3RIF5zpST5kBOz4YIsGkvoEJKKqm6MVFSF6m
dWGvc1/rizKtQYmwG56SEx20qz8fHGBbBDazUNahvqfNy1DlJGiAsSFLSn2WU6GrDTP6ewOWWXV7
mb2rn2VrTv8eR0myQce6wa/2PoAtT05j1qwLnObGixm2EJadlzBriGGYb4d4OssafBbdpPXuwtFI
tRk9oE6SKqO8Tx3ahs4eiSOY3H80G8mvu3IJOlWPd0JupKVWQE2Sl3ZSntYAEQ+M8S+yNgNUFJIw
hQlV/53lG2juHapfKNOJ53YNnO7K7peIeMZPaIb/7vByKl05nw+ynGQbsTf8leN94IgrI3LgKVOz
CqTVVT2KDvblyNoAEXSJp5eNPirKDZ8uDH6zi7WwX3ZxEDBbzxNZexfPp3LeLfay78KnOaYjCGBI
jH4FFyvnuppTBhZ0fT2+JIfWAqL49+85jeQn7htbSx8WDp6NbsODKUps7xD4n4cgF9OE98Y+PL1W
t1kaWbY21iZXKGNFajsTS/PO21W7nrAFJAsk6pd+8tP6/B+oLUqbr7a3A402zxBNYn5oSZZ+y2L8
Z8OdX5UzPn8pieTdVs3F2YcKTDE5tjZbbfU9d/d0cpK3eA1K3EtG780kLKgQCqtUi0wgNR5kR0d2
c4IiA6KYHoftuyJb9FsooI809D7cKEPG9g+gFIv7SKMx+5ZPIRCMrRSgIDFzyhOlKaSfdOrtl3eK
iFQlvMZ0YA1N9RSE7N/3VGbs9rOnY4gUfxCaLYLdwB4/qlY/RSjHvxbdWoRmsLumqEItyxlwEpZN
tHbOr4tZ/0UrQz08h2U+flzHLkW7ke2llLUWBc+uRUETP7RjjSQxRCaQFg17bPhJhvEcVGeboojS
NyxM5/4/IzDsrKhfnDh0euLWn0WDsS8XMgFQ9MPakHhAnds0uBQ925T5cVAFl7B6T6xQLopCHrXu
3gJphlAj9m5/uPCARX0chBnxY1EmkhcS7ZvOEpejZkIQD7yy750IoMfzogRYQM2rJZ0iFfYd9ZtY
9MN9qiKwgXu65/l9hSIwpoXyW7SzB1FiEZh+Xz8g+pYzjO36EqQFt2fHKP2T7fJ9V/PJHzylvRj1
h/vf1KM+7BrKPM/Eb3PnZATHX9xD+5peBjcjqkCPCeX7iRDWwbvUk0nqsEsedWxGsh2sC5YTh7m2
m5LUGUSYLfou1Ho9yYXP6tgTG4zJ54WllR8/uHuWO/uyOvV1CrNvUUVHV0roS4Z2d6pC91ggwpFw
q4pxyicAObxI7ItZCkZ2VWRDX6Jxd0QdwGZMXqAh7oqY1AIoz6UPxXA7/igdL0iwcdG9TdrTXqxv
//VFcK+uX0TfJSWCTO4Hg4ZxpvwO2Dbwf0OYxRglz3pqWDi03+EV/C2GA9oCbIQkjcp3Rm8/nqJ/
CIVlnaTjAC21xO09/N8uwMR52qfvGJBW+/y8SP6bOoHXLKiBEWQLse0owHVKXXCYU1IlALUkV12x
bVFu7apjlt8hAHrg27g/l8JN6v8oZ0vLo0PYnCZK1bbR71JpSmEsVgu6RXFzroKgy/RRE7D46iaE
rxLEbrCtZPze6BsM+2fU6ryCZ6MuPTVqU9NdU0OQUFzHpZA0obKeYJNgoi7c3tqQwSFfFMZTelWB
WykV65i6eUCpGU6BhPGgePdcDqJD0xxnjdMaU1B+wMKrIVlDoplBm04K8DEinKv2tV+m6FK0f+zn
hjY2laB8LUrJsRhM5VNUuTwsVNufx9inNu1dY/G9omy3sVsa/0pO6Bovm0jqqVQzsBKTgHTHFk6L
tSBohVv99I43FJ+j+Zi33Q64vLv1EI0w7wbWV6uSEgBkwm0Ar2LUIyui30puQ9afFde196z2VFxE
HRDF0ZZ1yqWzxDdfgFm8KHKJ2Kfjsr7EHsCUK4I5fX+UTb36JAwD6YpPsFEemPSVFkpsEWi/0Tv4
tOQWTyL6YzHoU9dQMAfByfgjsE4OBe3AcxyGbpr21hN9wFDd+NV/eoyGLcJsQdudLqv+Iz5zsuBO
RB++Ok7Q904zgzSUe2/cY5u0+59bUzZOWk+QiUbV97RFFcYYJ8jzT2RFgwODEC10pZrlj35GSpps
FMDtz6IpQcVTmkAc2gZinUUNB3tZ3OYBy9TySZEIe2tfztJT/ET6kyT8TapKLyVPRhU53TztmGr8
jXPPoZ8YbCidwnLTqh39XnwdZ3/OqhGRZTVjzJeb6K1Y21tno7npWZeLn0wEnZeoQsmnJIiHYrWs
4B4JhAHJ5jkh8+wUJwi3HmrX/3iISEGlEgpHCUs/tipbneh2Mj4LVoj9TZIfGkN5sKgsjZQ2ncO4
L3q/HATY8+c3ZEGIGUvS/wSCkbG+rXpjFOLBeMurUjOxt2fTKY4sMqt1scomaxM6pEbRsVesd/3U
kyr4poXkL/8eYE93nMxmFJuxsxez+f8lsHmYdKdcOKWd72L5E/ajgb37+ub8RIkm+kvYMy7O9Vlt
05LUm5JBCxI9zwWg90rXw5zTUmwCmmg1pVe7PYF+CKUgxS1ytSMZiZwReb1SyjMbanEIterVK0Pb
cbWNxW6x4ngKW79t1aKDJrpCcuJWBGZ5Zbhy0Fb0nXqIctCIQTLGTVHHw2cIUfVIdgvhDVdth65y
U78LNlD71iu4lFM/yga7Q8wYz4w4pgrcyb8FLHw784/pPulJZ9NvAxrvA6i0nMBYl7rfJ3f5bjA2
F41foCbBGpKOD3vBR8qcIkt55njgA5xpp4NHixa4r4T2JNsmIf/CNNH8IB4okdflp9lP8RdSbX/N
cLb0XNnThqUhWgJcb92GHz9hus0GDSPg4rPT8xUDToFWlqKRj6dl02yKscleKmCZqMN+3c/KTGpT
bzdFh0EYHQcMhdB5d0MAntG8P+9p2U1Gc01ZNYRlTPFMpNgtOfAB1k5iRK94h9phrNV+FfGEJFRx
2ND/8UsWHHCBgD4LUEkCUUGwAQW/7EvT22QPqszbVNbaDwtBNF3blE2mBwMpkb4xxPTE0Ax0bUDw
kvbLx5mRRRHAZDloncuyV1dohRQajL2wqSXS8c9cCDzz2nFDnvSJBNRrC4Ws5xRi2jZdPCrzkSOk
opqJBdfDItkmEu9i9Ymt6DlFGcwYiLo3OIh+oHiK3VjfNhj9zVLZSyZXIXBH+DG6zN4O7UCKDkGF
SRrF5PtKL7V7FOtjsfxbi+FnMf/ujxpk0TLXR4Z53VQeeFqIXmL3q/p1HCGvYppw8YXhyEouD12j
HqqNqftSFiy2YGjSojNY7gzdjbC3NQmuN9YTuHc5q7XYIKc6iXhUSxctqfl7gcSG4NSCgzzyGplr
n2EECprVkpBaJmF5pSN/jR2NueQb64XYh95j8/5hsgPKma6TtoTOLJiWyQfsUXIJLGBcAbfl+Cws
UOJYAAhCfmOvjQuUFDBB2S+/sbWAN1k6gK24u5hHsoICDx/63qog1WR+3E4IqzrIUYJcsyBEn+Ud
c8GP8n8rI+LI14u+Hhqg3bYqQdHPEiphL/YyzXsRYbHi+dEORZxKTuhvnzu0eFE1CQS8ege73rHf
WOHplc+0Z/L2LuNv+/HTyB/R48KNZ6+yzeSujHUBD9/URlZD/aQsreO6Mz0c/VhUnfa6ghMpWjcp
XmGqkt1NNgzZF6wLIA/+ty/NN+FR7+BR9Rwyl5zQTn4INuNfRrnZJi+AuwmW1j+Bnnb2Cqo9KYTU
NtQCMwML+Yzfrm313NOpoOv5yAb45HZuXKlVxunnHWrS9veimAcKWbOsXtOd2gX0ls5cFb+PR19a
0Ug6tIYM395tTTiHG4p+ZSUchKGKzMqqO2Y5/Y/LQbDpB3AS16kdXcRBTuYt7wL8r6AaaOFLXtzM
YC1R45B+E30E8hx95XxwQi9VIyG9hkIsTIJRfWsnjULBNIoiAaRDHd3uFERIKlquzNsaHtlSdRxi
3E4ELRzuw/FHc3SKdAGg3Z9eqPWC9zY5r6222Ah7ptWVLBkC3+DInFq+FCeRU67ktSwv/mu5FoBR
rXv+EjjLqEcMD8Sq8LUgEvwrGZyPyb9GNiL5TvDQL2CJGL1LvbOxTxt7g2iT5ghGdnbRVby4wvlB
zmRmxUuPt7DhKSSQeSpmWCNW5YK2Uf+9+3gME6yah+ELlft5lVWDCNP0LkCjGiRIvcVxDd2GxI7W
W+HkzqGmRS1q1vCCEfB9y+FiSrBwIfcw5LAfZPTScbhEDoTKIw0P06sg4Jr7QfQSMXYmKLw0ACua
uUTGMfrnVhZcLeHsshDQlaGPYaGcf9W4GNw76T8hNeIHcavSIde30LdyKTbKReluReZfUjwTXM6U
yc4flM7ENAYfb/CKTIqKAYP7xjw/fRCE9C5VuoLNboK3ddrkpVBJemKaUMtW0kWTfZJiPexcPB80
7SrqfUl5p8XL+LktGPxdx1HXvlOOZ1rQVDg/b438dyDTe6vXy23QT5kl8NG5pvNrr1Z5QtM7nqeH
aSRNNqBkOmnrKprEenxlcY08KtW7IDgpoFKA/F70H2KSCb3Ko+PVq366XaQkL8WGE3Q6DaY4R3pt
mibysUbsUqK+O0s8YJfYsDwidbGyr9vEgQeqBoxkA1veuuiutWHigxpjT51NvHlGQcubTws4s2a2
d4NWBYAHvAwkb+CqCuNu0oR1V5cGgmSAeewyBdaHvQrEbGPm+sWdQQ8f1Cd4MEz6wlaw9CJyNlOc
ogbv4uTAX5Q22HxbOk9tSVujKoBnPXYj/W8bH0ZBlMmKXuK0ZgNlhqLlEC0Lg43EcGSZ9YkWZQpt
pBcX6D/M5nuAJdPxAzwtVmUc0YyIs5uSnGTU3DWmbAdeldwjAyWY/bZhpyzNEkNyrANsXfPY4muO
EHhc8MMbYJs8ePoCAhw3Mi8GqM+2weTkZg1RI3IVfkuKCMuXpcleIS+wwjUtmJLsgTr+Gn6/jxUK
fvPXjn3ykK6I/JGlPUfDs/Utu/ajSBfsAE21Xn2JHJIJSA19l8FVkT+nvbzafoV3ZtKJXR0ei5Qy
NPNY7FeH8BXd0L0B0UjsnHtNEN7DvjWEkCstqNmx/fgZqSwWMk3eUD93/zNpW9qYtNrB8kbNZACW
vpdCYTsP7lUrvF1nYyQo/LqSWEShojynm4yiQgeihwzjd5ZiNKgnwrD+EqZGtRb6FiHUroXFb6WL
IC6ZjMVdQ0QiWUAN0sQW1Nntaou43jvhxloUCje6hEKxdJ7JrFG+HrLv+PvdZAjLD6yu3TG1a8Sp
1l2vHV9Y/VCjU4Bdm8x0Z5bLCpJdCrB5oSWtYWcDglSLqBjW6A08r5lkgp2wMDMqYaNSNGdka0xo
rWFTaNuunCRJ1Lf63r/0odz0I5EqSFYiwujssfsQ0FnzIVpdkyafqg7uGmnrxNGfRYESXn3G9Thb
HPIXV9DhWHz5VBQ/OUTWX6b0cq0xR/sV+XuSbz+pNO6WhV6rRJiwQ0brY4mmW7ij1R4OvicVgMbH
m4zxE3kej9fSpz1w5DmtJ07knjSTGPQsxxt0eHJoNPz3//IXoeL8RoaskFZkCig723dn/qWWEbtC
HeLQ9ct44WIz1SZUY82n+U79cluLUK3v69RHbPVWihWM4t23TetBlqayXtnSFvejlj/wKzMj7dem
TpmWQBTvzWjBRTaDHuHyDMCiZ5LxCSBriooF+XznA6YhHkjeGNbh8k0vuks2qL3mjlNkJBG4x0DD
Eh5nP1vyk5ee4aVs0UGBg9BcXwwNKsdA//Xsyap4B/R9IzQCs5jstgoKqWByIVrkCwmgBM/rOGyG
YJlWHGmiRy1WgFuIpM3Th7lPqjShs/cSHHStKWTsh9J/8ZGioIRtxxl8KgA5UHc6LxyNhC1+YXB1
y0ukHoB7gsWDXE6LuM5mL2a91pXA+UX9UOV9yKfEs4fuDSCXjORM2rvdkQQqYyUfSY3AM2J3eX82
B5y7F1eqira9z6pzaq7LO3m65avqnE7+wQgGq8psoZXoupsZ3fXcz2TFP8Ylt87xCVEnAbanLFh9
MuX9UlWI9Qe0PFnRY1XbNxkucoyLFgefdgL1fl2YXrNwj020tDVZyycHx9ZPHmg/ye5/YsQtEY0H
bvxEcuWRggldUN6ary/N0pvZUqd9oZ0Ksr7mQBbpH0rr1AyHu/IBnWqSUYCG0fcHmJKhHtQfm4rQ
h/6EV31K1u7hF7yZy24MN3XZPkNGRJ8A9e9fpd7seYNWTFqvPnkt2oZrxykCJq+eY6+5To9Qg7uY
m2Lx8G9Aha23JZ5c12NHrXrDTP6Rms8S+sokg27+emYv0RaF8c5TvoMQ7tFSpKvQbxuNiu/dxGsA
3UDyw1pTlIlBed0/UFwTyHCACtgUfLlrS1wGOgECcOpjCyfSditeOg4cNeGSmTfzlNn3mt0QENwz
iX+BTZ89nR/N+0bqOvqK52TWGkBO26MxAr6BPKoikcnKrVd99r9B0UAfTOih/eoihZ2VXOgA9NNc
z4yd3P3rFU3CYEtTO5n25bE5m6wwi4fYXP6ZEzBbXlk2vuXpPhRTTKJ1go20rWHijPQMAY37xj6Z
DsK4Qgo4ADpcrJhVnvAIBACKSxfmh3cUTeBWqKxZFlIaEeBVPEQG48nyJz8H0zpxBAlJljUA2VT4
ePy7XDQ9zg951QB/PXYeT880rzlmgP7IEA8V6zDuG51xnPCPgLisMCozFN1AXojyZw36Oac2FFBK
dQ+tXVcVZYTmO58/tQiAwwYHL3kbE02hjf13xx36A09BIAjJrfnEWCDr2olM1c8sRBgQ1wXhCYe9
jsZlAVh5kL5gQ6Watm+TEHry/4QMG+ZIuVZY9l2Q+BKoZVYmJ3KMWnKIMJjt4E9UHaKF0tUG3RuH
EtRjoPx3caNVKI6DS8ySOkIZRVG+cBJNh9CRn0a6RBIfUt4yqOrKH9XCgzEKRua35FKFo3P4Upp1
boxvtXAYJyTFreqNqmeBfdXXeF6vtjJUUaWxcg8FkBwL99yQlZjWzGho7u0BkH2GjAbI8fTnz8xr
C96ywsYSWtq/GY8jFCrQz+KSVL0POjv7+lGmQi/AoKJtKcsGxQe6VA7VB9w0N2E7VXFVzNqiXN2X
qLYZbaUK0dK1Sccc877kFM3G0GhLeVIFeCNu0mCohvK6zGn73NGHmMUPCVXR9AVbuhPFHiOkNoUf
5Kn6m33kwrXBK+T/DDK7YOXkIvAJ7K3+aIkZzVscOKF0Jalj7x8uOruvb0zJHPOBwAfvhSaU8Jbu
ZF60jh9jTdy28sV7jRvnYcwsugyvgSNz7ch/JSSeJQvTbi1U2lCLwVywlTul0nk6Q7fG4Ig1oYt1
LM5RksGAOAZXKkso1wlVKStYL4wgyEnjaLR4gNQMOEIiG6xtj/MwLg1DKxAawmaBOud6t9vh5nN0
I5YW6He4L8g5NUMnyI+ZZgdNEiniH5n2HSU9sjVXvX2oiwRmmrDhdBtffeAkPPCCbCgrp5Y4sFGU
Ru10z1dqLphbnVCt1ugOMllDIikzv5jAkAUs8saXtm3CTxtInvGZBZouoSWDu9nNIblWANHOeMUG
ZXYIfAXu/sBChJb/MW63Hq40d3t99gAIVfMsvhXcwmNjADtuMYRtNlXBFeTwVmsBhJFTlu6N/sLW
gYihLIBHdwB1GaXwAXirr8yl1wNLodE0zPP1Dt3L1rMVbZKtyP0J5j+1N+f+XZg1Gw5jg27yQktG
MDB6B5PBEMmH1SvL8CJKySPvWYcpTyhsz/+1depUDBLpEKclrmszDxOIdR5OmKtbs939Hzcmb8CJ
dwMB8WgwqrecB11YfdxoCiFf3qGjF6D5wPoPdER2s8arhmmWiGEphEDk20TDMcVwHYcViX32GBAG
GucwC0UZBPlEdryQ/lcb4FtP5atZkb9QhsOLB4R56GC/ZrnVGfq3ISAD+5krspp2tFs/PtY79I9X
z83vB5ayHcPUHWk18ya5OAqreS24M2X2c4H4bUBjkCCVNgdUmVRFNS4isF/jY+ruRKznzdzx7pbm
vFClINBxAAjtz/oK9bzJJcgnro6OQDwip5c99zKcB/Dxfh4OqwndcZXUEH19k0QDLTs+GJ786lQg
ZqhqNOTrOfchdqib2kq7hLk+n/prioAkkHijtGPNQDu4uV4dLfQ4HbtKLI7s/dLuJjzWybXYcJb3
LjD6YANQXmDpbwD4r7PXB2GO6B0wrFO71lRooZzYLZsDVhjx9BLgki54785Pq6lxQbmx5kpEuvEN
7NvfQ+nF+8WphO6nDAvi6juW2ul2r1y1wym4H7fHyhYY2y1+nMd5h+kYCyQp5HId1YI7zZh3dclo
wj/WgJA6u8jpgEMxneElC7lcVfIU/RnCHK1BRVN0/MYXyqof5mXDUVr9MNHoQrChVo8rpGBROw3+
sPwDf0OnAuHwiu5bEaFmTg3D8Uq8mfmDii6zuqe9g98R1LxKOMiklIPiK3TOxDoCfzC0moCVSxDU
4c2c+6XF61ft3vnv41vq2fj8dJNqX1nNQKAGnD1ZSVFYiIzoiK+vxw+QC0m2RV0CashHLO6BL+yk
t9y50se8Z3ipbrTxDBE4aX9KDJvVrJLLuT5ZVygfRomdLYGOCPauje1e/LFmtsKnjhfYA3wNPMiU
ALy+Nj/JREjTm34NgavOC479GrfNfVocSuub4NU6nNB2a0Zt+xPS2Sggs1Tw0QgkVpf4uZGKSgk6
HXYFY0Mmp++qaAWLN37GS8nva2qGTwxTw4k9DwfdcSq4iXUv/cCSLgT8pVcLq8FMcAX5fxN0mmLC
Sm5+6WyW+Fi5SKnlIc8BXL7R/DUcflx5zBN0mnTaMcfA1WVzOtrCjNvvQKyHcrYlqXo0t6aAhz1A
gOIqd5DcjOIEgYLTOMPUTvVJkNTjC/qhS3KB0oJrIe3tcokqIEZNPUX/Q7KzIi3JOhShevvERokV
kxzLH8H3cbvR7TZYA2SDDEjr+zvfALCqxJnnoSUQbgCBvopyWcD9PJXeSPw+HQ3lKcL5qFN9FUfT
UCXo1bEm6XlFWmf6gvjYb4XyKjSca0fwUecN7t4bdAOiawad/hphib15hIKuls8vkDqMgaxnx4JG
ZfSTn/AMht0bcaU7SfSN08x15uKrAG1sXM+Y5AW4X5lxaV3xrnkH6okB+5WksMgyLm8GK5Du7vWI
2LPj/0rCSV4GoZ4RZH966ztVEpzppfCwjpXw3GJo99dsGgvbq3MgTyLn2T4/228MNyeie7clkb06
XmuTtLMpt+ts90dyHcpl01EIdwJpqTy5XZYEQ5OkiKrXqFGpVnwE5PEs4zVGHgB24yKqC/D/rWZz
0MO6x8hGz5irk8nSX1FmPUa8gRlbPdDspEQojZN+CasnOJJSobJJT7Ix1dk4al2UL3BOCvERVsdp
ibpjFVehIjnXeL0h0ipiaNQp2qkZmf+T4FwT91c25hWvyf1pCH8k8MlXZtMMqIYGp72S8AI92ZOV
9ynv7WVaefYqqt100YskBEM0ISg71e+PWURDj2i7ipl84/HZa995P2EAMUNfblLlmbHjp4ShwRX5
0W7xzW1ISbdGwqAgNvdXSPapBJuLTt3kuefa6YHCnsCoKRsVEssIVZbLTOXpoKEcLjOvIGW3bEDI
NYon+1IuXzVMVCcSFDdKfqSKqCteC5LBdhq42Su/0hcms0ZK1TRw2vfflheGuWWqzUJjoBK/I5+k
YCUyuKn6pmUOopOGm7HvMXrESe6VBQ+VUG5pV2xGybjTjTozVGPjI09HkHzrcXAGCu/bkHn9hwy+
p3H0UrAs9u9FnMPkl2lKxgZ1kaK0QJ/PVc8nVdgmQoaCX1v3mClHkFagyA5bo2pxKeJxWPtviXg9
Lr2Eo7ek3Ya3ZXNdi1MupAf7CRq2pTAHTEIRZWegvcg5KWac/VDL3bdDsL7s5oDEEI/A9MauUdN9
N2wpwnSbNMlJS11YQXJ13eiPtUp9f2GahPEr0DVrVmcgRLFlaF2V3jpXO6qbxqu3tiZlAVWg2qCL
jYAbNmv1fEZGCIA3I8lmro3C74gNbtj5Cy5VlNe1/m0hEBwX4kiPVw4wI4ZyDXiYWTAP1XU9URDR
T4ljz5cxEWqlJxx6OFB+d6o0bUjU/cc9cOheKuo+oe1eE6Q0vz3xUqUvriBenXnG2r9eEYMcKuZE
aziZItbLu/jVpVBuZIdW+AkQriXORM2pYu7qiSh+b4aSpBpbPwbnCpTWL5FPsZ2VfTLR2QDNnDCb
qZa1McCn2SYfB+0sqPYNSBvbaj0pN3jAM6TlJU2A7p9AhZla+n6afQKyN7zQiJ/PMbW0EHsf70iV
o3YYxqu5GRo8YVmPTbPGJxWGc91VhrjgzhfHDMjakmUxtvbbg+FORmgL8OWfKt20HjKrSn8XW2lZ
Rw0Mh50HRQxBJ9Ioz71+/xti5cDyCC5PGOzJXCQCsHXHkPx2cqC7m3N1B3DcMKoJiHInVMGU4MJZ
7A6SAVlWKnqKH+wB5vhUGfq7/E4Q6E/X39qh3bzdzAtQiQKXJlU8LQyZVMdkaFb2Mg/0jHFtEF/X
yACFFh5bg7QGj9ABoPDQMqPg1IXrcoXmS3PnnHIDV9XBVmPCfuEngs9eW+BbmKklGuPCvs+AUeRV
+D59Mcp34mMDay+drW35CZ6gggQ4ne11eS1h85+NW2guz2W6/oHVf8e3PN4hAFyWqPv0bKhK+XXU
eFlItnBlqRxMLsM00ngjDXDjq8QC2+p/t5OzbL1LCTn2eYbIy71JqQNoJ6fLOBFFUi0r2ajOJ/5u
Xqw4gsHNHPmra+hHGAoWJO5bgAhAORP1WH+qBJuy5dR6kJhVe7lerCfYMzr2tp1G7xExLnNja3R7
yzQqL8RD2nCgjy2QH6wH+3Jrqt/Oes7TycfzVmHO1MoMLqaomRHp2ypVbWLtsjoD6N+9D9X09HuG
TUSiiGx6DRD/dKQwTRmLp3bhU2aOH1uVWrVyJuLL8br+afHaAkY3iXq6t20V51hptS5AWMnQbfR0
rzt36bF8tDZ8Lc4sjQlQYLoeKHqF11F9PenRiEvQrcRwzO3poMaPmQhMliMZH1EoZvU98FLQLca7
w3dwFjjwIIC1iuZOd0lSYJ1V0ZX/8enN/17YsgDt2ZFBDNoHNEXCYLtOXFIzj9liChHf9234Q8Iy
0uo7CLufhul66XfPYjGPzP7fkNQ3YWKlGtFHnlpbeXwIMCMUqNOV8vQ4SEEroTTS7a/HGvHMv+zU
9MJ7llGBE9M/eLrd74yV695t6YvmYFv1si0MAGXgb39uNn3l44vss4wPDrdkyXx5XNxlKfY1A3Q7
e8AplpF0V1/NSHJwRLb4GHtw0iByPngM5y5zoOA6S9u5zRg8I8BJG1qeLvNvpgW5ftPuRsaOnGOH
375Z8PII69M+OI0/TnWXshclhk1Cpq94htzqBA8uNfWNkn8Tnmi2t2zHiJhMgMGPRtJRKC8Hx/LI
TIv+Hx2MzKsTPMClfGYN2ByJtnOvIiKJ8bBu1neiuYP5zfc55UjYwoytM/KluOGbEpcSU1D0+Yqo
9RRQr+G44RXXAKUdeYAC8zYu1wUBfBa/Zvk2rwkATe1OtMfL1EpAlzwxMVYAsZyX9YMLkMzJ5RMP
oCY1u/a58xEngHCsS60RoM0USMvVJsLfoYGkMqLgdRL2Dpy0FCvG0Nm6Nhz55iZ/jzaS3shh166I
hbP8+l7E0JS7ti/sq9Neb7jRSXev1R3YoEkRdTtzWQ5uJjcToO53B4AM3Uu8bDR/+NFXJVlzsjVQ
ttVNJ8sfHOPukpGcrLiRAHKvjtZWUEuylj9eAywsM7ibNdNnPsHZdugaV/xVFMNwByamYfjio/MX
fE3hjdewloQnPqjq6X4dARHMugbZGrkRcbKijjp5O9WfVR2GsEVua81+PFijaa/EA8E1hGTYh1x/
QCffHOaZaRAZEty+6t6TVmv5fNgEX63CGbOfCBBXIWFQ/wJXZ5RkDcv+CyJY3GRCkBZRpij7f+W8
Jv9l8fr/iDqjaYGqzKBJNhRuS3v//Z91DTF/rsWgtY69qqT7/BiCaIdLa+ZQqjgeJETTbwKKtrxM
DZ1Hjabuz3MQKbA04w2ry4wGQeX5CSwnX5csrLj4BVkqYUqf0mc3qWLTuiyQILRhlwbbztLvPpKk
3Hc0BSTKffhZ001tmZpJnnj0zd9RB+8nAQTs3eVmKFiaxov0/IZYFB7ZjnNVAwCJpYF2yI2RHJwA
36T3CiPd5Anqbu3NoCP6D+Ew46hLTN/NeX7bMEgKcUiDsklsA4ZWCXq9t/qF/cKx2Z6Bv9Nm93TX
vbmNW9+TM8NrPdkkY1w10AFrLjPPvHI0l0vig3iRdL1SrxaEGLe/n+c1vu4Wdoi2kqX5A59BdtsW
Y0SrsDco2biHRQgVn/CYXMzgmEiQei01x5ghxjsd3C+PWPOCBbN0XnXio2Zn7ZZKSk0T8FTiXrw8
SVP2+84RUibo36/bfapuDFKT+otOehs0v2F5vc1iIQmcLLQviiMtksAobQSZaB3P0jYjJFzCqfKT
6R+ju+9W58Rr5bUW5hze9GzvteotGHOCJ/G0jEC2D5tZCZjkyCzPMQ1JfuKHK0U7M9u7CEWn/gpl
yR6swqnSMKJ2m9b66zG1mt7yuDldIdTOS3mp0sxlOQarmt9k3MLSP06juijins1JLiTJECKAW/qI
ITJTJQCt+gUdBShI5zyJSR4u6H3NakYsPaKE62NLtqUVV0OCK8QL73YJ/cKTXBQUJ9fPvP7STvUc
InkN101+4TqDbch7uNO9KdAbkmTqPSoUWXsoBTH1eIgA7ZX5T/6I8xzFOy9MaiswQoqOF5fLwVxG
kqvVNfYwRaiz05TclpYFDaOFKiht9dYcfeUyWjfWuTKaqWA0wjLkmRfnC5SkSHdCtC8X7+VA3tOR
+M7tF7y+wTCtTVQN/XaQu8HcitrDkW0TDezJtf/520bbO2LiWU5LlYlnv/ZlkIIV0O1rClRvj3Bg
p0f4hbTH7rOwucED5di7FHKupP40VkGYVqo63v3DteU5jE1Qn3phDqW+5nQhJrdcvUkdt073ZIQ+
zF0OzV+IH5gPurX/kZn/Fl/Kvctt3zFyHItiSRLKDKP021UmRVTYnRSjBJpLjbg+h/eCT+NYd1SR
fCxWHK5G3Oe2AQLynfqW9XfpopJlk9GSdWLMEx+0yqREhkA7ZywqngqEC8IL/tGDYYEU/+vqjBEa
O/NGuNKj01OBfLZLuzZEHsZcqL80NuqPrw5Mbp5E5YDMlsYTl3/EuSEOoeUjmMyDxuygEz1cPlrl
6MxhxhHKWTABNWsIrirBINAar6HLWQ/UUEAv7t8WfZtmjKnkPPz0Pb284OvbX9alc9xIYuYllRNk
IIjKrfGV6QZWHi0NfQWV5cUtgXNRJnI3rryVGmxecM9+jOmIaURRHzA0mTvHZNXsmYmYujWnqUnG
gTXKowIopLaXvB3XtFSf5eUWGN0oAZKslvNPKhmo/Ocyqk2NnJa/lNI4z+M2MOksVCOX5ZJNykhi
FZNVfFXUgmJOObnyNAP8hgYirUBzgoDhdVdl3CnIYNHOW3j+Dx2m7yL3koaW0RvSkASmUeTz/sqW
hKoDUS20Vm12XB1PtkvoiryLaixYnXWEFgYLwi8+J3ZX60qIhTGL8NsgX6H2gpazeD94aHr7Zojr
abOrnNo7qyUzIfkHjeB1p47phX5MfxaCsGqW/XoQdoBzeqlz8qtoGAHtTdb+3+xh6XrXFs5lgp+z
5GwmPaCVn9D5KJgRL5d1dw8KeLdAs1iJY5kelVkPYn3s+7bOPxQ5yndGGQcwBomFa6o6T0XsZ57A
ex+wMF3xn3NSFrnCl3lAsW1GihvUqVdeXpwUKXfrtlczDsilWk/6gSEh5svTG6tY4hulADYR/463
hq+dSSG/tD3yFogToEXQnNQ4b8m/sa82SpfH5kogbOTyVzsx5zr2esfOQFeNJJ++eYXqgBHNmJXv
A0PE1ujL7l5ciwZcV9AtvVR6YHDkI00+2KdISwzmwZpT+91uDAzK04IgZ9a4i5/iUc99Y/DFRd7N
Ys+i+Hisbq/7ZOZuUhZ7yjj57jgo5ojjI6G7KnXiG34tQfuI+XbXvR+EOkmXprAFmzxjVTdzUBTD
TBtEBNIz9LFWE50cMZiCxQb5BS+c7imCGuKtvAu84MMAkpMzqv912ZIKm5Y4whn2BrSR+HgZqCFs
ahx4xlKVylwwzZeSRHpC6nncuSRphOSGPnCNgSOQ7BqyziQy3/FEObbBUWqyBdT6ID0bjTPAm0if
6ExrW0pSu+ye5LK3o9Q4/gIDsO2bp+HFn+AIZCXktW8Ga0tQvcKNZjlAonWtKze/A3bdobb+pSIP
EIaXfNqi9YYe3QnePdJtIb5lFm6Yg9B2j3aa3/MhWXC6GlFIDiIuWdTFC6WCbxEhlsTcG5LJrHLf
lKqONpujeTQ4DsTrd+8E13w1GJCXjDz4K8HH4Dt19B2y/POsIoSF1kzY5JODkR428hT6Zau9VcZ9
vSqz2jpbUqEJ7QRMv09tUBdmRCaouHjlg/kJLaNsJEAx3B5y1P9zHP5Y4htvwhT0NaAwcngyZMGc
qCeFUQw0soJhpaY60bddOwIZsbY3/dvGZL5LKgwtenxdOdZGdAIqz/Vp8ic3XFBr5KCfdh18HLc1
JxeIozElHAB+NgwK4fdUYySr9U0OibdXkdQzvRh5d+B3gs/oFbRc8Ea98u2/yDijSql7wsQ7+ntN
tndplcAXEcIeLmzZxclGwdTGHshazY4Tm393hP6WBfj+S/3iusCtk7FSTA/qGsH3QHC835bvXuSa
f8Se2hZM6pJVe2bPCKEWfOJ0tFw87tXrXtOptHsoqh77vuQ3pzWrJ2Ze2XovdG7utdzc/K0ZjeGy
nfMzp922Vyx7HURani1WjVUsOrtKtuvTtJHhISAc/CD28Pm3co1epm9nQ5AwTp2RvIeEo8Tl5LbJ
s3OiVfPWx/ebqUuUS4wdYZc+qrYDeVz01KjzSjkYm4VtbnTbnL9tdrohAgFjuusNIqJ/1uGD3l3m
PYpDd13bclYxOouSELzGoResRyumOy68qR9RV4Q60+bw4kIG49zWZylv3QiCt5YjALOqjBi6udRy
Z9+cAcCu+ooKBZDgbObNYeHObeer7E8qiMkIhRdoMuA4jnA34gNLTEcX2A2yE0v7hn+7bL6s+Fi+
1qaQf6vkQTZm6Hp/F9nrarUVEW/443vxBDXS2C8KXBnBQiArVZkT+p+3o9O7WWv+aiTGANgtwy40
OkCvx1k9lQ2KKgBUR1KmK0kQAug8rLujQ+w+rkJMg0zikljsgfZg9559zaLS/ucg77pmbNnEB3jS
DJTINAp7LXIKslLNwqdDrzLV5lPfwYb3dtZ7JfRomGECy2eQpwY2GBSXqtrLGS6V3h4Vq4Qpz3RV
o1zObvpZ61tE2zXISk5aabNdXUlCtn5LfMqUcTjzkSD5etYemxrQzd7XwY7Ym00nT/cbrDWoC3+c
C7qd/+CHzsWqGvOkxVuHwpVJlW9uR8ruGbv5VHPifSV9zov/LTXj52BVpAiOJ19fOsG6CAhnP8vV
vk5+Oysbu/lzCnfOb+22lHMVnBU8rZrpyn3kmyz73E0YDjRu7/+sC91hpYxFa8OhwpL4vOINFa3/
DRqkFhJjJ9FHoEqoMZGy7x7Mov7bs2gCEGBZEefXKC+aiMqGJ5UyFBI9DXDQugWaDS1Nkzrv3nvk
E+ZEIIwpjaHc+J5wIQmS5GvKhDuy0S7Fzia0yq5lTWc6iCBzh6vMu3xVystEu1cl71J96X5QfbI+
/472WsVx6X9KvX6HyoEgQKcj/uTk/LQ5tMpKF0ErbsIHkUr+67xY2WCor1Ws4e3l9c2EczvzZQ6e
8LFjYYOXvsIMl2pe1yZ3xkQJlCYhupavb/Ditd6fQtFUsB9Q4JZNCXPqyW/pFbwUWIm1w7mQUKwY
B/DPfkZGxicVCGOIo2I66P+Vq9zPEhigV8b53MXvOnGs+BUpm6hq5WvSt9CosI9sUcKEPhY1ZaD2
TStL+TZsiy2v98377YrG1lFl3IVOVYBc5w7D58jGjguNRhUK2tBeb908Jh/g6mm2ylVgmE58c7mJ
hJAwkngdFW+G7QHV1bmydE+gwJmHD/6+n7Tdthl2bDZhNtnUJKTE2g7ixQEBACHVQg8v2gLcAWJZ
ScJQH7pUmX5oxTBZc/lFz3Ya5a0d1O+eTjMZNymLB0rXtyjYQ6w7FSrZGLZMDo0CJBb4HA1yjbpE
xRGPsby47HfqKId/u3qBtW1o46f9P3PSHrKMOzDiZdeqzT1HjTTFYPGGiMXUNNHCYfsvEciPz1OW
W8910xr/Gn75oTWZ68CmNubCL0SDeazOh/k5WFgdb3l70urPTmt2KN8g5hOqBQvjKSHBVNh2nAiL
XHr1BpMT1qR6T/Zc6En5NmV8ZWs8yC+0GoBWqI+vI8KnhPm9E/dzRzrR9Wl4LCm1s4/KHdwvvAxT
Sh74/s9fVgSBFgUbZ8f9/EGOt4++6x279iWAsiFpV6Kv0Z4GGTQMwr8KfUO0+7/GL9gKRXk4tWYN
m8tDN75QPX/RH+s+mj4XtqXyXmE86sEkFmHbTybIjDPN5yNU2CWDh+yUxDT0oUpSsX9GYKBpH/7B
X3s6k0gllxMRKfqeJck6w3NzCNXq/9nmmzSN2DKsXADmj8W1IlGvTYYPiTN4du/PtIwVBVP3Q5Go
ECPS5+DPFdg24l9tanuvS4PDtrHw4dP1bGXDYh/rVsKhTsrL1ajgR2BcuE2deSzDTowaPqgZHRsG
w+CsRr+r5fVPMVEAXqCH1BmvWysOzREkMHzLdCWZa4pCGTbyvQO/34Q8KmPuw6gMTir7sn72z62n
4cJHJ0FPto+16eXUyt0iAgl4B49iGIkkLbtEBVeyRzuOsyLpcQDJxYOANY0TNq9U4yKTwd2XsnBo
KcvKFhBkh2+CWU3WKR+Vxu7esXOzsNGgEWwApfAOZCma5Jor3k87Mmo/jAChSunJl2NK7QEsReOw
OZ9L0JO/zaqDC7eyrvggWR3JH/15YCgDtXgKZB0oKEerwoilLMpJHSo+QkgNzWFeXvp5Rh1z0UPE
TObY32f0mE6x4CcMAHWfSEeZbXOF2uALV5yGmQcu0CzHNnJ1GaxvZTvhgM/7K6d4KZvcDIlKzuC7
Djr2SnuxtZuGNUojhPiuyQhPSF4BOMJTBhS6H2ildsvPnwowySFp0MihosP3QeMVmub26wOwEiwa
+D8HU4BouqDzlHC7XV7K9jbs4TWVuUyMpIdq2fb/oyn5A2EyJpGrFv4rkGDmlNBsdviNiXEONL5v
MEcKmdmvg1iGC4jf3LeGANWhD74o+5lzwu8acGl86XOLZ2o+yT0BNc+C+ggHABfzt8iTkQHUm9m5
Who2C42X1FLsXov/WTTpS1cSqVUNKmA99fOQmHAIgSOTerVX404N+fHzxmYxAmwnMS4BWsEn0YpW
lhrZyVL95JPn/WViRRaQxCxsZXqAnb5ZhnHkP+3JsaDbq9gyIwsMbFkncVtse4ljf2hYUbwrT1eR
LfSTIJTeLCrBoxbQpvCDWnRJXBrzIpr/7tStAeS3ZBc+Rl7XiX/taPWDyrnT2vcQ2Zz4DUDWeq0P
AQ4FdMTEyX9HGCuunRCw8NqS7HSr9uXHCaJxYIkLuXnLHb9VcPeBBNa/szS6a50xcrS7Y06F6rpj
HOO1HZVkTVxlPkgck6Q5USYjVdAjX2DmASMnf4xYdhpkuH5bBp3Uownm74RG7hF30RRrxWbjlW+/
8X0/9ARpTHdgeWtaMtA+aXfgbJ3ewTpZ++A32dYxZTjKl/p/5h9vCf9YccKCaZrHcjdb9Y1gcOLO
BH96pcjYKV1NliTIQhKOphl9tUm7tk1thnJqJfeTIhTW2j3KJLzFf8SpEFGBweIbUT1KaibZjiLk
LUmGmZUQSzZsmuuJ4OJ0okAsRk6SKEPEXtoBsP9knio7kCBk7BPU5SO6Xise40mKLzDk/Gdox0Oh
O1KBCVPV0K/cd+mHlwCXagefvd9Wr70YIDRCY5bgeK+KTu/VeDXCqsW1y7Lzmv91ljJjwHCHtma1
n2CswNsp+MHshxdEeYO6nNSUd2zjuuJEc1EPZYiKqQdxsYtUUg/1ca+bJx2BDot0JqZm2l3w+ane
sOaD2oGn/AwSvyCPlEf2av13EjlGhiyOYv9+ROCkBlwopYbkBLtzsU27WMnYMJtScz2RGx995tNL
eL7a3WrHB4pWsJpLXwcgwzjSQwSZQdmQW1BjH0LSWKoSp3V6SfiITU/XN9hIBqGe1y2vS5GFiQKg
DFJpIO2+ITVKX+597F2ndpvkv8HKULkq79oWxSFqTvmJLdHC1X/Lzu5WDGoFXiISw6aVw1iGwfdm
cMWGKXkNpSCCdrCEkCXaa7I8ASs768tAXfwldmzmVWuxceCG1eEnHeBfiqajYmQziFcXqI1IAZpQ
FQ3LfXPrcWib6h1FboG0sF9YhyyKApyctAxdzt6xQiOsqqyrf8F8dx1ReZQ4j2WXMHkgSAnEcBSL
1IIHG3zD9Gp7DTeRn2ODExbNfK19c2WImnGm/m15BSt7OSXPMTH2XxGp2IZngwu8VXKxKZbsxtBL
9OlxHKito9Li1ERJHJ39d+HLoqqmHibUjJcGfSMlNNfodsRlR+tU6xV/6R6rowBOC+jLm7nDatso
ZUiQP5OnjnsK+XbSZTkvJlcUsGSYdnOrt3bVMafKsnKwmY2plndJpvr/085DxmSowcnDrHRXCpk1
HU17XpvM1xAZOqQfZnif1GAzDFerjkQaOUzWthAhnNx0wF8csvhKO4Tk7KoLjTcVR3RRjrJocAP7
hhv6x3WUgNMh11rs5BCM0A9pvwR4kGvjhletQeZLeoGbPNiNNm1HhDGYooCD18x8UOd3ziECi8pz
XoBXHqipDUBbKyxqZChhlbf2lJNbu5lnt2w9yi2XkW8nwCCBTpLKGpEN8JOVMbCKxXpJvhBirRIm
1xfQ9plJI5Bi6jdIcTUQYimfIZuheezzQ03iJRGI40pF5QmJB2yoENiMzxd0G0S1F3swIfqpROhN
XWDKe/zb/P4z0BWxAXEDwYkYYyXJQCSv1aJunLlNYr3Qu7HqEC49/wAOd7xdGvG5wtJL+CttN0T0
jRRsA7jq3Y7u5BSYS/lDYTJ6BIxVLO0r1ltB0zO+MY2FgIuoFUgpY8NM1/1Y0nadmCVmyz8HKaog
jxWWgv7NyM3w7jlujGb7lsmfs4jX+Qzl8GbGCXmH1o+QQy/MZwHhTht7xpZd/xPzJ5pqAzi7dR64
q7GxSQkCJMCRs86pUz7C517VTqnEtZUiEChDIG1yj0BpNhbYwwwPNvD6FLsGeHRfhT8lzTPyadTD
Y4SrqCRARRPdbdFvYFGP5i1Yt5lrPcDMk1ni7AlgrZhdCprzegFJEAydnzlqK29Srw0sHPN0KcUt
ij4Na8/s/ZijSpe4KJnqOkafgbPnVHHH4yWrpW4LgEGpF4rOq5GPTq27OwP5MdmKqJCLMNyQj8dc
0zYPaEBMRtDRTIhBYiSttmFSHVNlLQJdyRjlpUYsphztJDpn/Cfl7QLhz8SuvD75GBepl+uBFQ0w
RlaS6BlZApUI7SkuzSmJ9k3dwAODlifnQ7JVVvGWCvc6DXXOoo1sA0BaEqAUMID0ppmje1aNei76
TC4XwcJlltsUMirfQ75Txty6w9zDICauSNDOFfsw8vlbcZtJa+l66nVJVDlBhywdELw8BtplnBlR
WN0TlATNR2fGg1dQgFt/xXrwF9GXM8+hKcxLHDqEzeQV3qtzkB47PnZb/SGLGJKOUs2SD4ifUQXo
GxZXv1OSSSoPV6shVSedtqSEvmqFiUCY8dutMUi9r1h+r9PtAEOM3OF422W6sDXeIm0wFGryhzqq
s6CGFuFolWOxGdV5hBbgcbQg/TfwaBU5HEgMJoiKT+q8bhXe7v6NTVRuLvQYA7L8r83ARXmVMK4A
lAPJFY10zfIrpwYh+IXSQShKkfVLt3opNP3MXN0HWbQBkqOkLIIxRDkhUxvfKpYsW9WLtFuOh+Zg
KVy1zIn9eU+aBUQdhUiPWR8ulMe+4nGLodMNPC32Owx2p9r+LM+fCBe8j2pAYYi0EfVEK7YqKm2G
CsIScT1RFQAM3UPZr2rkHuOTvGrT9Ly6kAycttlfglLLv+4rmYbvAP49LMNqa9Tex+kDCrO8PS1t
L3q8TyvVPDygHDfuV/fFQad2sVt//Je2fYTumK+FNL1OY1tDqBTaKwKWaMVdGYArfP/XQQ4OrxTu
vHCAIsFIuk3WfsXS0LyuOA1gPEOz8AhaokSjPEw7aQDxigDnA+xiA1OY38NUMi3i3WglHbiePoni
yuC1apXriqxrutfMeg8Azsd7fsz9OpVkzkWxxDdgYUB4nOebrf4Sh10U7GySA56UEKkErSaLy+eQ
0mTjXnIwAEI2ym3SvdiK0CRBIQW6JsHG1HLp/ypgqxJRVLVtL+vCODINUu2Fy2B9l1W7efRB+V31
kQE0h+z8RIsaoa2+JKoRXQiO1CrBT0RzRLDG1ajd9M3qPl8bkzg5WqYScm5sOG6JOv/uHicMsZUw
5kyIsMDUqqEbSW5J4OYK0JTbbcLOOEpqOQ+iUYte3qZEZ7Rl2sFyhCOksoImsMbtLWe6m03F6TLp
7bSs/uPoEXT3TW2sNH+S8Dx6oCuuqVlo2qemCdmTcejpPJmw1dVSpgmVJS9ASb8TqTYn3Jk+qD3P
UaIdy4VeodxIydJQM5FF4jtKuamoXLfjJ9sw3ljC0YFz8YiYWLYZH5c4htlN3HNzDrBFN8jpH361
QiWw8TJC4qDcTVs8jyCIi/26HhIkDIR901SJWaz2RxvFPXbcUa/Vowe57MA11hq0wtln9nZ8fo9W
r4QfUm62ks5uj2ecANAHQJJ9ciNJp215HwC2bjChu3+M1aw7P5t3Ll0Q1P30UCgh9k6nm2gEtZko
OFf5IqMPSfwEjmUhpx66e+DlhlEpoNOD78oeScDTR4qmxZ7s3OKfbPWH76CgcWZ7oyKe2ZTWs4Lx
TOPq39bBI+NaeBshjbcx0nzSYCNwJu3WN4wQ4G3q7bBnViBvaiFWUBPY0KPxGEyBaFK5uXqzlj0w
JxHfnVUKDUUZw1U20dlOnLoeiSjj94mK8F86GeCz+BzIK0ytDlPbaT489vApnCpYgImCPO4c0pD/
EWpLull5Yn2uZFAbCw6pOoVTzNfD67agqFEvqHpXPv/rLGBCUgsUzRLyHOw7DHeW77MTGuBUpXQP
2DIbLFpjVWqJsLzUqLNI7G1naeLFWOIRIuDayUw2DxhX/AQKkT6T/xOP/BPu/C4i0VL0llcUg+AQ
VPTRl5unHeMiRJfjn+4eO7JbSQ6PQm053Oi3CG29xF0Jp/A4fD+ag+OGhsrr2lNz+0MMdOgsY2mF
XN9MVbOucIbqX5U6mZSKTEuio25hGVjGV8lhZ+e7IR6jSxQVDS1rG5ea0V4I+rBDHoPJOuHHyyJ0
aHDsAvmH5/XiECod0Yncz4ULKqs4n2CsNz1tGCaZiiiVJg0flcKceltU55RRJ4d3eOTSTxEJh79t
8tl0EtzN1D09ecCB6EjOqujh6Gd+qM5caL6nQDDwR59BzyVCcSU0KrYyWaa5uekFkZxPQ9/ao9iw
qEo7ePsuu8ACB5bhnTLq62b/3Xh/oRVHWcYMChqILTO41RpTNNIhrvmQ3ask0KTTHfk2D/eAJGs4
Iw/73REjDvt4A6VBPnwXAc2n6x3YBDJUWC54BvQ2FS5K2zcni8/sBQv93/hy0BqyU/7hPcwR7ctS
yjESvnNaAdWWEt7OedRlL2Dn4zdy6nj/rn49BaD/DDQE02mv7FEUhi0j4hfzBEpCVW/fb9ST8v/w
LcPYLqPDwc29IE6hyEKSIWcklWFuMeVyt09DLRyNZu97Wdrl3ah6sWK+COsBhsr4zghHuWF1S32O
+RnlpWxL6yx/xE9iLTVBp6X6PGSU010VrI9Ei5VRWExue2h4E+GG2B1LGNGUnAfsHRBl9iJf+EFk
g9Bz+IxkEPNddKFjeZcPRG3mj6ZTlaJie26n1QKhPJXqR1mJeqVbPiAL2G56WCzMUw3BcPoQLqBz
PPYWHK/DoLfdKZ5bKNbX6rWGOSFAAPM/4bXaIVh6+O4H4B36ZZQhmnbJXb1nZaTjNx7xY89U2zMn
VMRDbyUq4k9uu227L/fIxtwSGm4fuhc1cqDVAhyGO5GL3LBOdBIUwVXrfA88z4xxNA9tpfocft+V
I1sQ5q3hCq8kxsHBo6PBDGsh5VVlfWJz5SNpWGHM3aNUfptOgwDtrv9HqAEYORb78tCwMl0M2ytE
WUR35uW1W29unFwHLbWc/lsvRoX3QnWBDMCqmAEoseD9fwOcYcVrfKb2Nv/6ezkgxe/t9Xbj6u8g
Ec+hmSnLNxhAgMAFSsGbLfIsaBMZLTqRRhKV10cAEkvVrkmiFXcZxpE7HMPRA7GACiKr5DLMSPB0
1UC0s+SJ1HcpOiqxySCNjgfr43MD6G/jpzvngYcdkXT7jGyRJ2AiqYQhzx253OibYJqhj1x8J4Ds
2V54ZNeaLCJb71WPwr/FWMUvPpo7iUU3tIXO9yK+gcsbQ8MzbyYkFggc/G+3Zd2VsmWDmDMa9sw2
NLNw4h3A430EJoGAGgUJAAoFslbxh/tNnuviFtdb3ntgFgzLiXB97fXoT8K7uTSVC4f6WXOyNQul
rXpVkNgxCL49PhmioHznAq+0apGij6mKh3DJykfyR+yuEGKMcKCyvcz4TAHHwixFWvs249xdncda
qvH3xya+0KCAlegiif8XsqbPVlkHpBBfJ2n4RgD8Rz8mBH07suxyf1QzyBW26anLTUopEttLBapR
UeFPAQ2kE0/qA0cTYDYMdI3I6z33gSTHniZLRSN3JxIu+axoCoAi8crClTfxGHUVF9Mp7tMjRXl4
6b0yIeddnjdo6nAg4jbCkxyOX1P/hLj8LXWokBE0VeGBL4XdJRg9mGSsVLJUQC8hK0R6e0yEXhYm
oEu/8YC9DxjBG1iojUFR6fypUBs7fznEbEOuj7gNLa3RxAANTYM8xEyd+wxg+s9V10up6H9YAD4O
gtq6Y4vPPqJR/vRVITU4vIYnGwZysSRievTiHlxG8zZdWb0NnDOMOHVLHjad8m3YGk3ry9kTsERq
sATVQBwWmmir0HcM7adXDofWw7EJJ3ezmE0rOajpCuGJDYmoYymzR9DomAjN9ChUf8H9xFUN1WaA
KCpHChWw61eJmxffV+FY6vQGsAFrprwQYy/WaHNLaUvKSx4O6TSTSeBMQhabXD0HSR3x2N19wLI1
FJqjF3in3c/m+xDg9wa4zAWNsQDF8cDHPLtJjU7GyOlaHeG/EbnjK5a4TG9k7ek74xVGCLzIdswe
3+WGCChgtYJL4RLcYzHs7ym+0y3X9v7Cm5KQUCLlvPoAjyKXY86jwoqt/eK0ltcgiEgs/vktiJ3f
6JdZ+gwsUh2rD5aaENtN3L1+MJkaEMeGYPHO4iJXF4k+MifnHN2pHxCr4V51K2eWn+FRSTlMlSO6
bwhM6pxFPaOAqUW/7NtLi6IqLGhKffZSxyD4b3IIoFrWna7E0GcZeLNaYnMUSDDZC/70ir4+SnJj
V4JPEqeJ7LTPxvIfrXEJJ0Ai06zrU+y61d5vz+1I9mkvOYbwfjr9PjZjcnfTV7tmBKeu+SIXNRJY
7zRO3uu9k8cxEppW3biAmEfmdxe4w0qk1nQay269Re4sLT7y4bZPajb+nVreAPD4/TlGhEMrVFKk
7DWNJ+XjhXfEJSTMTzRrADveVzOSMlli8R7RDGG8tort1YfE+Xl18Q2eLQxQOXE/DQJ5DzxsEecx
FeuMV7Bw6SlXDwQjUK9rN5cz2qYvTIt1U72wK7p7ncX7D53KaAhZp2ZrCrIXvlm/uI/QDNnfHf5o
piT42ahBy6eTzsPp0ToOHlcxbsuqRq16+C33B/JZT9NVH2ro+AKnR6S+jaCAyAiGH1Vm1FPkRnOw
UlpM/vzhzMiglGbr/NeiH/x2wn8Rmxm/WZnomwmVz+QXsjx7vRax3SwDqg0hlT2LBmrZHYHTIu0X
7xARNoM9Y+OTlo+VScNF7QU0JEiy+65MMdSUEbGx3mXlS9NK0TRsooY5H6djvmP6OhIFY6xLXGTV
aZDv6N0f02kj9Ip5gLm0fEvBUEgjZ/2Ir2o4KJ+x1Pbl4sKdP+PpU+FwccZWxXHR6kGHRkfXVZMT
1A6iykxSN4NsG/HYr0mfM9BYtaWDCoHkn4KYRtmxZ0nP58+J7yJNU/6tfjWKlmVspp8+v+Ne1sTs
j3JCuh496lyHVoXrYxpeJF+fy1BwJoJAEpjZZz6lorTdbuVxwIcA4CR4LgFRV37YBO4H7Bty2Kso
/9XoBaU1StbuZY9I2bXUOiT0ZmEupAqzbCncOnTIBV/TDw2o/Anud1prGr20tCRpRZvog/I8YYH2
QUxOAwnBJtWh2fgNaxW5YjPAR7Cl0EVBT1IbdHhQxI7iVoDnJigwZlAJA2HOusIhCBOKV8klIKu8
PgTqQFDg7ISWZdhr+0VuRUAXLOVv14qD5oTscQJAfClLDtyx74eT1lmnh1anJT+VRmPfPPepCAQz
+TPrDW20798n5xfWzLDD15tp+IjWlz2gK/bFMrUFFG8Idls8dVpntNudWqX27WFXse04bptQP34q
PdTN3hubsx56FzHZBxtjnQs8dKLzSbylHQijb+HlKglmguvXcMqjE77B5/Uz9yglQ9SD3TZ7miH2
cw7wvpui7p0T7Bw8FcrwOt4C+05haGojQ9uRGpLbMQuywWT+sxpOihHfN9O1mZGlWCp1IVzSQL2D
7IuSPZUjDUO83tWow+nzht0/rIVEwnCbMVBaebmbZI2BL7ofGb1BuS5evFBkb5/rjmwsfDCYuOtv
1MnIzNAw28pXVPu0B7Y+ujy/dKNTeyi5c8DROMVaZQhRHmkhVAksOgn8AEtiLI1oB8oMZa05Gy87
XcyEdc/+UAG2Xm9do8P3EfrpaRiconJj5RVaLu5KWZlO7B4kWKH/rPMVnfz/4kaIk2UR90ZgMyBl
lI2CPwA2Keqi/20VuwbFKsohShbTkWFMvjA2Nx06MElpMAUt4QZhh1cz7bsHttu7paCAZ5h33kiL
iNwQ4GbVzHGKwgBI7zQfw9v2qscsXJ1w1ybBjzgbV3LBZYIpJ0yIhGhKsgFDr7SQhhouHPEZwuOH
IHfFkMdWhJ3Ecd0iFfIaE2M+4pgkKWLfrHa09Dx/9gfkgcrJp7HUe6ka1G5hkQZLKnJu4zanCu9Y
79ADUH9+JgQI7F2QDeVo4ELzcRGiNq46GxoCMFX9CqWJ2Y43O+n35mM0AhXe+QbrsUz4c/cShlo0
rRwZb7TDVuntI122NoLMJkUDGVnCECOvCyYV8pKyRS8W/f2BJKoxdqBbXDzIZZmPstWDnpwTMKEt
S/pk6RHrgrx93SXmKNo4oTs8XplTIj9cjgKEjfCB0qig32sr8QB9nuAsTeYNJUodHup9o1W01W0d
TlQSfxeNIVUY3BRBA4B+LnBT9sr3XJ5M3LAqyLsWNZ2mXXEO3hLhL0Qx7D1g3P8rhyr1KS3QOAZ6
7k3XSjvChYVquuER/Wy1NmQZ5xfFYVkl7GvhrdmZGR1IpVPKym7sqc8F7kyck2E5eLE9fMJYGDfq
ne4rWuHpoCn/U4WQRiAjsELtT42+9VKl9MB0CPIyMIqJtpwvXYpur6/WtACcD/aRovrSIncWSBgB
n/JMVhjF/ic6501a/dROB4k4sMowrW2reosVnwWMlaytkih4z9CvNddevxM+j0GOqmsFe6mxT/7N
8gYcCFfb9ToPZSByJM4C8drejiJS8e1YH9INKnx2971nJ/IDJcrGH0ZmkUemoi704PD/U/0X0Pzg
5WsQYX06BAftGbvKonL8MSTtDnzApmg4XXcbz2+I/hCQUsusg9w1Kdq+JvVbLhYbuveU6P0PZYQN
cmZWQefKz6+XXlhhNbpOJ0XOclrjH0c34X2ZgoKtWZ8+XZvyaQt4UJS5x5rSS+Q1XlJiuztBdYwy
Q2gFYJmFSjnGeLKsOQtxqIefVTx9v4QuxhetHBGyuG0UZxrKykex64b23x09HBU1J6ZzyOQmwT2K
NKTGNzcYUHCtrAnCBFMarOXTBhOKRpeXsN4K1LpUq4bX7+Uoycb3Pax7B9Crx7f4XuHJ9F1vKu98
7ROo7EDGrt1TrlFMhe9sH7NTZB75sK+OSiNtAShGK5GaJfXAy03fSlANj1bc6O2equt+38lwKSNZ
wob2cCB2CXAHigR/akzf+zJkAYSlxtVKGlqYdIqwrN4u253nQKlE5Y9+eC/UmdNd48TT1UK2l5ML
e5NEt87NvexePfazxG6UtuwGxsQj2vqoPWmPhQ4DdIgunLXcpk0l8fecOrdJd2unrrsV3medZUdh
2zYZCO5YdIMpoZTWZn2g6GgpuEaRcmSwvaSL6rOmI7SvroEWzw7nsnngq/UFZD5DLsjCLnuMXe9c
9hFg++9PwlyKgD+QDG1ysLA8/ZrGBbcS/IGMESn/yq6Hf9Zfa6VNo87er/y/Ag9bXfqyr0SIe4ll
qIHOYvX+o8YneeKLWFfwugqQdZ56NubwLxU+82T+/Qnr7zK+T0Z5A1aN7NKL4aaJIPhEBz+5s03c
A9mDxcTk4FXHsECnGx5HwTsNLrfH79X0vUOeCctw8ekZsFIaC24hPjsME3ggBZ15GjvrcdGDrhCo
X+b0FacmQhy1rX8PWiroDcnddSCAzqL+A5pICeIN4/js+UvZoOopz+VytKDAVVXcGvveZG3WNrZ8
fRTaLhEunzpsZcPNF4y2ISxzdIm3U+z20RjMaRovcE6adyglsKJVazFvr5kCCrPwEutKGEJ4Fd1/
T6V+/eQ5g+rCLBm/mYeEJ38fXeMbYFs/FbM4Bheaaxpzdy6wUZsIU6o1IWcbqvt4YGJYLyYC5v1C
V8COasMS9Xt1OtpVw7dwZERHtZeFRPewgqXZFNrKbC5y0VcVlOW0UNEU8j8MctxkF8Yhnt0oNax7
nK6BDjrHRoZGXeG0qxv/LCOMkf6tsx8mNiaB1z6vJHwOlQ7xKCL9UzWG2EBPT/69qNvmFiy7Zbfp
x/QGnQesreGUmL8dU5H/IARfB6HAz0sppULokt+IQuxB2+ljPgwoJy0yTuUYxpwnDaHFfNNIAV97
Skd+UayKTNK3MQeMOTIckmiiAj/IJk8XBBF1iB+WJj4X93BzNy6rTSrKKkocZ1itwH58VZOXD69e
wr6cemNU+y+Jyu9X/IphzbkJ1RNldK95tpx01cS/xGeltODfgGf4WD3cD6zLHr6e9ra76pGI+qwL
3HQBzUgZIFJbHC4KYmI45aDCWbbdPRnjaLHkPHyvSsizjZod1M/8cRfn7ImiyuvwaLgyeDKSfBEh
7wDVHS6jYIC7WCgeLkEGVvWE7BTcKcRQ87zLmHb28MqyBaD4cxmTy5BZd0F7bAjCPBNOJfx9w1cq
HzzF9Bdr4EInwWAIpgtKZDWbpX3G3RpLaQR9/jvrD50IRXUm2CDy9Af8vn2ITYCSGsr7Pat7xv1p
idB4dO5qPtcj0XAJG9inzFTLCfcKrEJ7vJxhTIpapkppp7P7FCy58OljB/LxFFbR+weTMR1HxPmp
E//dX8+ecVZiT++0CRwWD0RUDskisOuHiJT27T6Oyq4y77CfWjxtnsEwbMBQ0kFAtUQJnsuxYQMm
XYc7iRy1hIN1ps7X47V9zoHmgNMj2rTNiMTSRINLgWVXem0Xf9vrCrD/I9K6BnDlQHIkGSyxmO4F
ZGBQxlH2g3gCspzpQ9nzds/fNqKaL2Pih3C2d51huqQjj4FrYihZoXilJlSdohEdvT6oLp6m8nVR
DFUUIdx8YZJhLifugszeK5tCZQE1M95eO7f073ozaTYslbfsdvExGmQWjU3zRs+m5XZEmH00Xnd+
Ef3NS0qIw+eeXGMWz8upd1ZtIzZ0GGN28kdjzhBnP+G65h6+GPW2eJltysNUf8J9xtV2IqYnkAzS
sfQkZQa2Sk+neqQ5y4+BxQsQEJ5wF/G6Ho9f4B8/80Th+hKClr1azFLKsKX4+RMfD8hvzd1OZOdq
BtBqz8aMZgiQY70NsJMcTbmPgNtCnm7Or0jXLnOvIn0ECYQrbQmruaZL2ZnKM4uZCXPCy20gyqsS
nZ2IbFB+GatgO83hNo+JhuxbKeLkmSCitJPXsIAyyfN7aCUEaW3LCsUPwI1t2+BX96CjQwMyIpAH
ykz7nDQ3mTTbPLtMIFTfDjBZs/8mR5zX3oOvDsug1/VFuGy9Z1gBIeXGr/pjKahZi67DYZ1lYsZ+
1gew9tHlYXrD0LhTjSjqevmimXU2yD34QE2A/H5BzwaO5roFxV2aWPMsGtGVbxDRbG7r68iQUNuL
qNr23F/NOuK/5PZ7E7NW7J40zW1SRd17IVe7u1QfF/nWutafMIgP4JONkpwSqHv5d3sew5kLVZki
5Ehc51fRuzi/bmvWryOPktDeNfQd9hKH85IqZRzkXodOJDZYpplPVyDlMrMPwctlE8XsRAbUwdQq
FGPaLYG7vyYHzYBYcqkqDgTZWF5JQyKs4ypFmDyYfmQ3xIGDd6qK6atigC3nDgeKsvXo37P5w5Ep
OAUYwb5jfuUxZWg7h1/EvEQIfmDorWmqKmqLqmuR5Ozz2u/1DGKcHK1YnU7gAx7y3bLtOSl/aEnu
KW8h6qsPTN0i8xfL1awg1iIL1x+uwfELVsMK1VXVrExpo5s3KcgoQ2d6Et5KeqS+yt+j1Ft0cld4
0cN1f41fjIGWkbCcyMnaQTQN6Cq6Pof8Fj3l0M7cQHSanaLZhYr07ATlI1UWq6v4uucRaJKcDpXh
CyEaCD0JeOPDmTikr48Z5cZM+rUNqxSHazsmJ7CGtpx3BkMvRmNDaEgYXlJfNB5mcK4dErYkMnXg
PfsuHVeEnRXjFREGE143y3r+AkJRVaXoPY8VRVSymNSGkdbTD3kxwfWmmzaxHGLQmRWuKWYAdIx7
gBWiAhMRBuWRkRPID9w591zDidD5DLkcXSNBebV8/nB82AHUVMFL9qNezYQ3hqs/q2cELJ6yiqPs
Dd2n7iPj0a6Bg7cgqStBNUgeXY9vZIiQGYQD9HpKSAYxJ6Nic5yPfAl/aDy6pEWCdjGv/CPcDPRE
MZWWKjGRPIdbxWUATOLaQLaS41QQVlPXOlzH/g7qy7KZxVFDtQ2Rx3NbnW1RfciI2DJ2XY941jZ4
b1RyY5UUN6LtGfky7jxqBp9CVZKvw5jjF0DJCiUJcvZRcnlLjnrAIiaJ/bbSYcgkT1ZUXlX5NFX7
jb6+wHPmus7IQ5Wm6TqXas/CDHfLKNp6JvXU7DmhzF8PLHE1sr33bsp9LdNrKbm3Z0EjmPi0vffa
VsMLUcnqKMqUB3cfAAIi+ZEg1KmY3eQ7S7wyAcOO9mFuqQNqeBQ53G+ebaER/DGMaeFECgPKJHZU
zeBjMXs3koPyPdFc+n3BG85MEb+OaX8hnaLJ2KYJGF0WrmYJOgq1wfx5SZ/VW1NKqxedParJ+Tap
/crrvbLnLc6wQEfGzdQb9v4d1NTVA3anHDn3DSEFwkgTHgxtX4wBNXzvjmMXlsTRjcaFhxntHRmK
NfKw6Q0MyI1Vva+aBXyJodxR/KNAzPZNd3eHkYdKmMEcMQjFr+xQIj1681ISfKPKrzW+/1OaAmDf
L3PMlN1cmoQjOZGDpKZcrQq1zCUVdhZnlv3SDTxG5puEWhLwXr/mSB4HwQqCQ8uzZuF+sdvHQreP
U+xC+Ze9ns2DqNGfl1QuXEUpOLrIl6+cHtW+SPMVPqPpH+vgYAlaxdEMdjzxZ/ahx/wOJpwFazQ9
fWkRAKMUztlO28y1mGEepsUo0w/Nsso1q7YCxoWH6QqFiOQDQ3B/2217umj+WEIJp/5QqS1XW7gs
Mn1VKsVlRN8j1LKCGfZO0FW/mdCft/4zwt+W7KSlozjjly4/a/zJ6lYb0kqriTOsiVZ/PjTjYcjB
eh02WfuJAWYb0sh3c26CdCwkls8LVZNNyAegMhSfP4vPou8IgofbMyy3ydybxJK4mrIvvVFN9SFT
qbqlqXXiHtuB2sXDOKzkmy/RR2x/sN5fsitQg52D1p3e3RmN6Q7ODlzui1Vt5RHNkU/3Jyyewsvf
Qn7Qm7V2ZPg3kcksr/cLs9ib08j9+hJPgnspO1O7JELTYhlmGGnHCZGRzlUCkYZDvxKVm5p2zSoA
VEvGdvNbESQWhvHBUspNhzmkwnS4Z44zlEChQOPTOh6KQ1SkyZeAWquyzdu9ZYV2r+74M5g7+oGj
6xlmgQPWzpO3/0uV7f664rmwwmrF8zD0FbVXRjkO8Y5aZdkGhiHXYvlbkymrAsZxv2Ab8qWyqSSe
aPlyGly7yG2jq+y3itylfkXhnhRPWbaYmAqrVVd/Fj8KOYYYhuglyLzxYU9/TJYUBJmieEu+++Rp
cLNjPgGl1OXgK+8Rw1w0vWaMl3HVMMCSp8+uIGr4eiq5Fzsx5J2UMtVyvfL1UaX3+07XWIAhFcjq
cschybaD/CYu/uRK
`protect end_protected
