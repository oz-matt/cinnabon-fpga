-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
NuMGcmMP+amgRQq8iBMLFYK/yAmcXsxozABWkW+k0+eGyQLpk/ZO/en5OnCUFJxys80z1hbFhDyR
Pe7Qu1LdzNIIlL7qWqczMgxECywc29CyDYBx1KmbP4CMAmXyguMtYkCGadBe+vexQRJWMe2iRJgM
JIfRPuXevJ7UWv7FKrZ1iDPE4MnTEw1opeKqaeRjYaOLsQB+8XLar4q0IM2D0nYkZ5hmdX8wlHOR
Ky3M446ospOhlf7qZkcBHWdx6/Z1lm+6RMiuDAL5JbIPE5CM6mHwdAVxex5KBEJW0ou6kKji/hUI
2HIB84CJptLo0bLOiJL8eUbAmzWbf2WgO3LO+A==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 18800)
`protect data_block
7NE5h3SxG6N1iBd8+BZ2C64ebbX+UfcUW0d3Dp13sVln4IG9cd7g4aZLDsOmYXhMQLvSGh8NBCUS
fn1Cbr1oEosCI72zTXWkywie7+iD204semzOV8wMXGX1VpL11vyJZ3p5mRLbi9QoNd5hIKEPyTDS
KFmeqG4R5qzR5r7e8H1MGjSkKKClJREichS2B+YO+IpbZy6U+5SRinykws+vCC/1jmVikrFJ9U9e
3fjfZldrwE7csnyf+s+QT+u0MZx3Plj3PusDaBv8BDJnbtP7DhgYpc7Zi4QBGsr0nMJ6bQJKaTVy
EnsS25fKGsayy1Oq2X5ZO8hrSNCJKnH18YxxkzXUnDd7PVMnQaHy6LKXF8SIrY/i2RfA877kL9ol
Qo7PAziBuSMG3OkfXfkjf7j2laSJPYAnROem5xTD+6Ob2CayLsEfuD50vSNOPnO2J/AcvNBi0+rV
tgxF5qGwOUyfjqaDM5wy6+8qzJ4TDdczL1Zg378r7tDvj6f0I9taN17QOgFMjGERUwN4y5eNDcnc
f4GZ8jv+yfjHfNz9zQiipd56yQLD2SIaXUU/3x3itAZWUugk/DsHFw3jOtpX3NFy6I0jJGdrXtZd
Nk8HedITD52IkoTUnmYpk2Iggi5w0ZO65eLRnjRpUgqKzh5ydwYTgqrRjKYCVWVQhPSIVkVh2lSM
AOyJlJkwTV/pd9RMGGhiGL5xoqxHWik48EgWVaiY4aJCtpcMAEB7CBWJS7M5qMCgk91FsfM3e/WC
oxXcoVA/mg1GISN77RZVybNgeJZExKkQeFpuOQTGfVqgoQdCKp/2ofsAwM/ily3qWTqS5r2xjXr1
n9BE2OserA4szYXaW8MZTSfOwUBp9j8KgGvQiqMoU94b2hNYCwUCUCmlWKSDvIBLQ8oue8mLSga+
h6jegiCuV0EdW9vkASc9NGfjCTbmxLjcqo/WdrFPJEJKgJjLyhGUTY+vclABeceACeoCKhZG/zXB
a8ezcbRJ0G2ZmgCRiT8Uvv3dvLXhpEQrT5LBWh4/fWi15FQPQhfHZ+eZJdc2toCv6Fayg4FCkUga
tgLcsbdHVne9S8Slfbs9/2rF1QMDyIERrXMgjxmdHNzKYhgy4qsKvrO7RvGD2CTlU1L85MBTvDHh
1qQl4Yk7SWI2yBweiuSvaPIBb5Zs26Y+ycfHYaj+4ZTjAsPR0YAi5aplIDLYiPSD/sqhxZI66i3r
r1wRf4rr1EmiPhL8U3BIWwTQTtHYxsrpu2xPCesUN2ieinQqWDk291VhRVPHs8xRbzc/DfhVwGg1
pxXl7tGR44cHDkQQxnKLdg0TF9to05UFD2iRHAwLeaGxr/TFTsKfXcyGrYonZ0+tS9cE2/BfLqQq
3HqEmVBuJA89eTnWovymT9Jn0IYNNd9CSNtTTowicsjEBoEqOEDXOCmaN0MxsvfeMfSCj8UhW8/k
z2BEAjGmn9Rkxu3TKPqqmIhjngVkncDNQD9dbHiiHSAOvnq9MZqtx1rk4sYxvfMHfrRArng64dC0
IdfpFWkIEkrbCx68iQ4fdI1V8jfjudBLOo3G4vUK2uERaHJ0XG6hKn5EKb0d+8iIhv7cQU8+YtjL
c7VAUiH0Zm/IWbvOqICmfdREIPuXmFNutLoHXWSlqT+Is6AwsFNBIj2F6c8RT+RZgi49BS39joeu
yxcJwD/2rdVV/7cwyKsTsQF8mFFHwtGZK6bCJX3/5QQ3sWWNi9Qopx8ORKdJw89tdxIpQMMzFcDJ
4o+/C+RR91NRKX37FoFf2if65dOJGyMBwJ/uetJr5uzOf0mYKg/QZS6xkPnDj4AE3RF+EqysSC3p
N4JPB+e/rQRbbC8p0mkfAFiRd1jXBB2mwNCezhJ09RoIXpLIcG/1a5/qpfMf4DRmH0lOCgFXAI1R
GofdbVRRKWKDMnbuwaRr69OsWoC6zuz3oLeVnSar5Ncp0yrcBXRs3kyqYbDSwdWS+eiHAfeTBO8t
DvG1NT5WeIyMz+Fjt69SRn2VrR6Za/9CHmwlaHR98XLEPtypHNH/ZUsb61t/PQj49dyv0x/eYdi8
EracGWNOfqMKjeQvXHtC501S54woyUQVQFfq7MuWOunRIQIaXYGD/n5mi6xVStC6gtyhclvLDUev
iY/+Xqh27x1aOnsojY48XGV8wkr6Y1vL+85QbFQXq4ymDaz5gVUye7LxChNjWuSjfqW9nPpQTEMv
rfwq8GqBgzx0h5Z8eV0DbyS468mg039WBoHu9CDI+C1dk2ZwdgijhvUruZIjjBh1GwQiEfaW1KDc
a0yy+qqrqCT9VenIKN106ULAJbrizpnJ9k0z7Y73IhjrkJD77kHnht5eqO1TToLSx8v7EGGtBsTL
NaiKUYRGbBAQymsJvciupcbLeslCjPwx9d6o1vG35hB8zHeQfTqpBFQNsihGoJVyRjLtUhkpQkLJ
gL4hsQ6ooS7l7EOzU3DTI0WzCfCQnGBGWtXhNBZEW595R0HZXuFlqecGsOOppt9nAEYzFIvqx4gz
sDEZO2mBukyVztBMRFZkc+/YaAVcU/gbWIRMnCcTYXn5jDiB6hU1hbC+OsEKUHtQEUmO1XwPFh7M
3JkWaSAXV1THmzpV2KNM0GYGTXhKjgPHDnPU7nhDenpZeTAdsN93hocrcoi3W/FryXKZ3WWasCLe
A4kq9FxrLn//OQThZ2R+qWxT/Uu6O4DONOARGA70gDDfFY5vxGD1qHIaNKmgzW2TMPGBa2t57bS4
X7g4zzRW4F0VcXfSAgGeJTP1bedeRxxJCmKAn019jUHFbAhSPDW786Sg9SHQWnw1SR5PfYiywH8h
Iyn5nPjm3B4h8+vldbyJb7IfUQOSmh5FOjnRc7C0Z+eoKNWr/zJUNzETiRVwuw4CWo/tKS738Y4N
N2/o8D3uFuFwtLOOhQJdAb5MxyE3O3DdGNxIUX+zlgXjXo6vQjbsyQ9GmdOrjTLNNBs1yRMztW+1
2O2kNo8du7fXtYBw7wMVpR9xLznDbbO5zBzPUFt7IO7pYeVcGfxYoFKbRIW1O2toZBH9n7YKH9nI
cbEBos0IRwO9HGSytM/dW6k3cOy6KBKHbKfMIj5Hd3Bz/FixC6CJ4zkpxJaFI5eijMFeiK/WcAnw
biz7xjDow7CJxa+JBHw5JRVs078h7PKpgtKgCsK9yPXXJL4UZWc8UlgjlJb1q+8WNwc81dUhj3li
Vc/AsOnzKBX+cpN8+VYVNHJkO1vUb9GWTw5QTIubbVp9FElGfeZgkkl++ygpwA9T6SHWYr0X50Ja
llpyPvtCimFBNLJwduYN3OlS8KVIbX+bXCjuylhH6hvI76vrPDKvtGL3SEw/z9cBLTiSI+CV7FZG
a92ZtdNyXwf/t/eSqHLRn4QfG3tey0H8XXk9lyVb7SlnSRRU40Gvh5sAQ4KVJf8h7L730oTMI8nm
2hP0zSH5vuwmBFcbvdHdyuTn9IlHtAvWerN6ifeQig5yrys0wSpBHum/kOZ/xucR0Z/u9aeq2TN9
UgUTw0MVT3ieP68n4QXU7bZcvemre7v223rbl6k2t3zYYUrpVlxVjZNTbVldRbsmyyniDejbO7/7
2V4qYmZly1Q5Rok5muzWMtjzBcnDgRkTYxGEHHmMmrI/BEhnIIAZJAulVbhRd/+CzablaJHZiG/M
zbNJ/BKpkvlrKf2cRwbnkzvZEXWI/cp1S33W5iCUa8RSre+HWPS7g0SmiOR8miEjUw/z1FZ6hgL+
cqwdJv2EONEEziUD1kZwOc1egX2qFacGzCT/rlnYoPB7seFylr2JltsNZFVfP9TFzH17x/Raxcm+
kD4F5ZYx6vbK0IT48Frb7zct8BMuYVYLQs4va28J8rjdVmIOuHSXbrrbJjQ3x0F7+TAoReWtmr6t
Ar6jfKPsPBu7IRB5+o3oR5Q4KjNjXf59x6a340EImnB6HKkeniZJE7UnSx9Fnztmuvw3NI99hBQl
fHBszMSAuRD38LU0qYsgYYgH3H3Yv1+UqbiAs3p5s1d312YAs15vzOUpOaPvUAAIQThmj6kUW8ua
/mwQdGu6lL+KfqPccFIT/yy2XRrBQsKLnSDdS8+8fbuJ+NP2Cfgn8v2fSOGzCdxoA+At7bPHZK6s
ulxqwRP8+4IFy69VRrDqPNC8LhDNIeydnIa58ZU0t8oMEGfevv1K+PgEwaXhFVgxpk8QuBe7cLhL
ADBd2/YCzLhIyKrzD4ZHBXgB1li3+Hg8S90hW7uXkTOyo3QSsDXttfJvkENNYWVT13ZuzaYqTkEE
8MksisUvwbBLvp0/xksLGPPdAJqzzlKF8+bMxLlQLjqkX9pZRHh+qzl0q0WrO/YFuGVgjwkY8K3Z
tJtyiAoTEmDlNTmYbIlOLFS8opujXPqMMR+jT540AgjrijVSNzNbpJ0J7WoQud1n0D3u4J4RfCXB
wITFNHiANJiLhwisreRh3/O+onrH9QBEUH62zWmWetQxZEOYz46GXiHQMa3YdpIs/b4AsDsyspPy
ByjHMTsQmCz1vHMNagwK5jh2TOILWwG3qr/T5ebPHrYDiTlm2yophsBZNCED3aHnnGs8gG549IMl
vNXadynORh+so99jdqykWMKvZTAmdNkiIPRhb4KjmRpqAPLLnctsdUnXVH0ooBwyRmJS92AkRJQc
CZJ6bLuge0PSlSAzCjOVMisFh4R5iAQsgQWzXEWbQN9Q7RpFtxsuEGmfeQzCduPe8pHuiECdca7k
s6tJ2hauknhwIsTAVv/Fq7Zf6KsFl2jqIJwKTineKpBQUJH7wCV1VENmamVN0+u33G1aFIOEu61q
eIfEBYpe36j0ELTxMdVV+C/Q4CBii44a4qawQ82ohor3KDpMBgDm0U0oA2O0wmZ9kKiUTfpws7hU
68Y8VI5p+vI3BlC62e3WI/gagRUvwxZgYSTEIMv8KFy2RRngecxAYNZmpWOL6EL1pZS1lHs2qNf6
ZryExizUt8R+cNhUIxdJ2riIsqWEHVaJmRPOX6BbZxPNm9oWKpWAYOdgjC26Ob1T3/xCvep2dzwj
7rCmE2IJbrqI6w3tPIcGcONDcgr94u1I3PRfiygkaB1Knuj6qFpDblxvBv9thVlMqQNLW2uj0lOl
uC6kIOLRA2Qnj+2W5xTe0MGzXAqiWj0N8OZsK1un7+h9C97xHHT0aVqTBZeqDl98X5L78wxWHkfs
wfc8iuTnTCW6Ti/514R+OUGlh/P6K9SHJ9r+GnIJab1EaoWcIr6pAl8nP79QJYT11YjX6JmzYel2
6cU5dijMxJMj5u8fIf4p8XbjGRXYWEjH9hPZBi33MVIxyvlQznk+7+//2LaOV6DrM8BtW6evckWC
HXlwRyDu3jLoJ3putGqepL6+aU2Red+rvQCVYQQfBSN4pA8S5Xk1d8kml8g5eXmT19V0fzPKeuJH
6fu8rodn7ZDoe4MuGAX1NFUes4k227Mf6IowzQ6BBNCQaa5JY7iq9fMp+FnKqrCbJPztbpXKWOfd
sriEpaXlZWyTX9dj2uTyvikk1pudrcpAU6Yr8bS50oWV7E+WJFdif1WfjYplOIxja81/4yjeDN2w
hTT10gjo+JPGK2/6wC5fMTn3tXE/yKzYJmulkwGE6qikgFbZ3joW7ztNxK30bZM/V76q4ZfrjsHI
os3usnGkr2hMvuqvY6RJ+hBGi5ZfATdIWU+Xsdwp76klLKpQymXCxy8PcBv3e/DNE8Jt2YfAhYKU
alyRB9kXg3ChzHzIlv6H1Or9BABUwl1v7ethBB+/jwTqWAJb0bYUYsfGZDzfs2x1+meDwHVfW8xZ
UdHgj0xD5Ge/5J6pXO06DJ3nyVv1l//HrXY8nTiMNzpxUi4nelEM3NtBRoWmGXNDGTSJQnjaxwsc
CYsYIQfEC6Ecym1gUO5plvMVORYkv1uYTMqie6BETPvsSxdaghCTjQmz6AdPZV4EJ/3XCKVFv1sd
04+8OoZOR5lhqlOUbBVkGr7WAio1JOFxicKGXUfljKtGLBAfLvKOZ6/ruH7n3sSY/EJsbWg1CIjr
eMdo9hqhG/LIrwdjJetAOMy0Lkun8kHYEGfWXZDmWv24HwyGDscwDPjYDyeO+5snlqADw5NYE6rg
Sb7CFaMXM9PinmbFRikQk/+iPk9SQfr+cJ3T4uoDpVoqrmNkx5pW6pZe2MbhwhbSVAlMQd5kfNtE
FXhrJHdNaO8jlfanWD9QQiYz9t1LvPTFAolLNwZZEIoTqSEOgLeszIXFo6zM6GsowtBjS/w1vKOy
DLt+KVVZ4Dw3W0P0g2qaqygTuqrXUoy7bj9ROK9XVELcTVsn8Y+StoheDUcPmdswxYVdDPjoXKsJ
f+jeAYDTTallOw4FCp1JGrUMijG4JOeHmdjezqd2GLp2KZ9yUouy/1HrL+4adcxsSviAqMeaJfiD
wRWYq1OzsWTH0dVBkOihg6XuU+r+2b+Pu7bKi4cD8Bkm30DLsJgLL9j7eORc14HoM/ezTn0CkmZ2
10c7titji7ic6DMHL2KbVxjoKOW+foXv8U+Z6xvJHjaMGoJbRx+FU5DMNxIQ8qNlFhpSPv7GBuUR
AEn7eF0JNmqbNNt0+y/ObQHY0w+oHVToPcLC7ojQ66vT1U7GwB+n4dAIKHj2kHxSIk9R9ag7TKaK
ikq/yqjQ7ZKiGVKDNKxsea9lk2n4nryjn/Tqnja/niHts5bhGW1MbqdGStexC1GPH4ZDY0ci16oA
cpX0Iq037h8XOvwY2c4/DhcClmX8dGBPPxs5qH6Nty1sOQKw049CwcQKEVAUzIv81kC0cwdPQ5tn
7gV3gDWA3Ya2MTa5e43QuSie2QVwqrjByDg+LS/TrkyqgeUz+hw05ekVTDkbOjYZ0Zybn3pOO5jx
7V5zn9lgg9BPSCLNH+fykrUIUPpgFyA5Ksq3MsRoJZGbtJAIl2Q6laykh+hhBeuu33b+vbuAyOtF
3HFvSghOpmpN6j4vgZ93PHZXup1SZYceKFnbvotI1nGu2yx/d6NCkUK0k9laN8zOUISrqhXd6+Bf
erH0bIe4J5r7EJRsA3S9t3+Lx+203c7d58Mkri4Cja+r0iEZyYhRafCG85YQiX99Ar0LQnIgUQME
/Z2EUkuZaVfGfuFlSYwilKLVGvxPa/tF+N6C8SjIZxOU19JHLjL1GC/OOslmeCjSPgLzXuN9WlNS
KR3A573Ek+qKDmnEDfzWQub+T1/ImhA87fkd23C9gEDOmJWurLXiDnQPsOwKGYV9euJvibhYxKbI
3piKWktY5UyUOs22GRFCzATPVqF0uB14JdOOk5t90ZDRE31ET36soMBRZsE3Ip0UvOzmSP1DEL7g
viQU2KmZlmLdNHB8GbTh9tGUw/QPFPQrX8D+F7Ru+t2U5RjV3JbaKiDhJ5Dz6atPjWuvXUsEjGSN
UAQK4MRIdusFprlq4QPNHvoXyhXeJb1IMTEK967A0TXeyKB0oF5n3KRboEnEBDdz2dh7QUCEo4ke
qhOT4nbpRb622g1ivYEQRziMx7hbvByYJxjsg2F58HZXsn1Jl+JnvB7NPzWhgIjQckSvDm0jooJp
s/rXR9/nzLrIpYrIkBQEliJpXDZfEb8uL9HIc5zD93QfM/0u0MQ0w3Z+X+7S4DJsiTsCAKGN0RAF
Rx84+ALW4GuboZutO1xaoic6Z1FZmstmeqNqcVdH+bbBghZ2s70J+ERvAzOh2XcKSQ47pnyxR05A
Us7aYb/Bc5TYp9gHR8FhS7WUcqmzqvr4t4yVfRxgDhjNgy8xqOrnQm0lLybk87xvQaOz1VHeFDwe
1T0oYEj7AFd3gaFLz6YcKmeADdjfA6EZHEFtfAJ/7+pLKnqijXIKhlJZCW1bP5NB/LCz8yBjk6rc
EcyjySXSiVd98LXtyqpstDXkwdqaw2y6kDiMPkdTzxDjssClyEMkqx/kGCAUxLP7ZW4QJPKCetHx
5DdqwthrEbsGXHW/ZxzSngALw+rnRDBnzyputsU1LaQJHacdYTg2bgOeUylbMRq8T2Fa9AM3nbcB
D6L4lC6ezezTabaVod5is21nn9JXvH7KxfuYhCn4Kd1Ond1K7Ra4cY2nWzXFYIesTZE8OBS4UR1m
oGyyMTmDO0pB9b8KgbpRzzCsCUf+aXDtDIflC3Ym5ej2GF8IYopeIMqwEJyCYwwSe/IZFolgcP1e
9X8wg2KZc5hI5+kO9nWPw702pPLEodqWsapOvZy4vpOiU2tKb3hWUjYfkmzkJHCMgAb8PED7Ga4Q
MbX1MZwLGZ38bgSH9395OfjlruMwJ0hOstCjxw7SayKQD+wRZ6znfvoIpc8bB0oywHE7HGWH0/+7
BEhD//FXXyR7CKucQ9bE7Nn1xHVaKt3067fJophYg9BpoVaCF3lwn1WvnFMGAz2ISWRqPNw/PAGt
gP3hVOE7NEyN6goBYe+TXwk5i5oykb8Om4lZo8koZwe/kjJ1Gina8VEz9w46f93hvCsqWBnN5yBI
dFoi7BJI3xL7qKdX40doJaDofDOe9bGpFiZyubKjYLxNjCnpzwA7e7Q9/9YeTBtd3axC2EIt6K07
1BEIW7SmYAyQR0BVAbDOBwPyOnif6TzArJUNtDft86wU5n+j7wCmihRoMLDlQfDb4oz/pYTthYYf
r4mhSHni77OO9psPNN0A7zahWBeFroHDzbpbynDEjPC46mJ5ERfpgbGrTnqDyqTBp3r7gzs/aC3I
IezVEJjuwOsA3ZOC5DOPiSsLHuLmPYEXK65ip2Pb2XsqqzSRB8BUrPLclV0GFyBo4t60Q2lf/ip3
omGyqTGGuU16nVECFFmeOAv0UadE6Fj7pl7ysaSICZT5/Xk6cS355m1pttrmRO3qcL3b+2dxbZ79
XWM2XdXfjqSR2kyjPN1IRqfJyAgtcl5lXIlQB/iVrHN60goYOy4+gUF18TndjGHqZvrvE9f0nHnm
7jWqjk1pZu5yTiFixPZ3srf2BuRGmnmtHj01YNg37U1agGUQUmpkdkpZ2lYo8+k5cgnI0DR6x+EE
ojnqobDt36+t95eyy9BrsfxSYR86iQZMOPJESgUidFXvwMtGdNeedVwdUNVstUXSmXW+63/iXANu
ANJ6otAICwXDMzXcLBE9eqsllFGEjxUgwDXEK+/2W9Y2qeLOnMd6kcY57SreST1qEVkALOPA+VBv
DbsBhXX+gcYuCopWcT5TZaLmevg6zJG5PxtURTLO7TgH0sKjf+8UvriEZiTw7SOuUpnxfsN4r2ZI
ITw9UwaQzsnt43H6JvQuYZKxz7SatM3NBJNe5XJ1Gv1mCMJFho35EpVw2qu2Cji1JvIaXejWXxWq
YLslXqxSXu4LVlRmpfGtOvbnXjdJ9pBdkYLGZFXMeEE53nbwN5otvdBaq28qCV+VL7gk1CB9B2Yh
FQvywGaM+pHGJQW0Jr4HPJy/javv+hQ+005bkoSuHk7mojQJMSBhm1sxSWlSA7jQ1mxXqnDlOmr0
xMctJiti2OV9HdHLSsPMiZr3cjWq5qAECwkrWA81mtxRD6Nm+2CvNMdb5MpV0QQ+w+fs210ihCTi
Bi0MdVuYwiWpdxMDAB9GbLT1jnhAHx+2ykd3B4WwxhVMmkKuJ6UDgBi9J+X31KFdCGPUzNKtDGbP
bHY+7vgSAYRlqiYf5/JzEne1Wdc7YRHeWfaWxiK3mEs1k53vH8DP7JFGBOpsmRgCWz9GkgKDIIeL
eg1iSFTgl9NE8SnPS4oP7h/cLTH8+AMEakrOm0v/Xs2C9IR613pufPqwraw8QyjGwmpG85xKbTRN
/yXXGNQFAnpJrqeC+t3Velgpy4TOyabB1JGZaJ6TsbvLz/slcmZNIO7T1pOoiAbPqgLcfmJCVz/d
HgTyzAEkY9vLt+Jq9fLwzhkTEhQVTReEYTLofpI1J4S76YUYTxEmChvQcL+K8VqT3IbjoP82MMuN
/Ra4uWqTHD7hAMcWb2OWppxzlbMu4aSqvxyVw/xJ0Zl0G9YTFOTqiMLMkQUTI3ALf4TC00L/O7MK
Yr6Y9kyB/gNouJ6p5HPOOWKnnpCHlOu6DOXsl6lV3uM4SF6KUC0fC4HSA/5eHX17bfQZAoTt4gYI
5XJdd+iybE5r4m1fdqXoPgMPbUvyeEoK6SW1gM9AOHIXwW5r2hntbRD84BdeFe7pny0Jb5ACxjQf
G1C54U1b2+iz5TFtyxWezTAYGSghrp7+/Dp/syW9RYFtoog50B+rx/mFS9O9Tq6jHglbIUAilYhB
uu37XWRHs1YLXL5wWKjIP8uV/CPANoZ3BSZ0E0l1l1tl+7TEL7q96TyK1y3uS3CW9nI1yqUdkKnT
7BX0n1oAsVJr6qDRk0GiJC4VAkRpzD2KMMweVGVxvJq5y9MOMYf0eS14koh659q+dQLvQU7p9ehi
xXeFD+AyNq90HG4lzWltq4nH9BM4xpaWHPMvb3L/cZG8+PifppjQtCDGSegHVTUWUkDJeDBOCYna
6cR+sJu9kqhgS1GfVx+U+NqB7S2qXkmBYVLCUBwBAKhBBrtJhFh2nzsa5qh5yCThcZ/7tclJ0qh1
D1Oe6qNjbbnTp6v7n91eKNIrxYQBkP+9Sa8SRmc1hF/o4WI8aoRiamOlVJwbPvsKMVxx77oXYL3t
G/GcVZ06adZdeKgFpkO7+dBDAVysPCna5elhYq/ycHUfBS4tjjJuum4LAdg68K2jHvnHt6ZV0P/N
0Aq/KHjIpDm/HLr/G8DxCMuQAtDNs/5t/v2sgVDNnbAVM3kSMNMupVdJ8pwNn+hU+EHqwjS4MKjo
Kdu1lI9wlhQfwXakQ7pKt+0ORHJGfsMzeDko9VbTFiNod4iXNhj1EoVnfChTcmM0gQkD1UxWXnGD
Gajjtu3UOI8YPRgsHlWGE8zR8WtQtwOQaZBz4HQsJMX/aRtmRPFYghUiMPglO6yduFfSVbrw9h0i
tqZ+aYC1LSptK4PpdYAdNOl11nFelyHV00ddJ0dWrSUd3XqW/XQAXdWKybq+bp7eAd2PHeXFpl0e
LbZa3j1wem/7+0PXcKYEdU+gVHW1Bc2Rt2VoWi/6AqW9B3ME1brmvc6CWtc/mzlMbhO7b+JCJ5+8
OmEK8loE6mJz6cNXAq9Br6SogWym8zNBR6HEQZkkfXk0gpoYaKTC0rOhDk1MJKJiln7Eqrd+Ad/D
MNbh7GmovCofSClEMd62+pgrS4qQrVjN1g2R0SmSwaY9C6zZENduo+iHE6h2icRSkO6rUusntQj9
rbWcxbRf+unjg2zD7TelNcq4blek9IqwT+M0X2uDzet427JqI/sVtahw9B2Zi719K9U+KLBupGh3
mERIQ+sFTC0M0/AV4nZD0x6jRBVbhQS3A+15n+O81a21H/B3VvLVnXJIG7wUoweqolVuB9QuSIJX
b/zdYfQ2n8Dlp3HEaARiWauvi/f/Vmpw7hn2qCxCqltFA2BLOY6fS06079otHoWblmPXINCpHsFh
3FxAq5QMW58MG6FqEZiadrtK67tPCJeVgIAF+VlGaYplF0Ig84su8TH7GxXw83are0wHA18hHkjP
ovKd+9izi92uupQJUphZM8HNCkEqCjkWur1Q2I4x2KzHo2A/gufS4c6YPh3ZduyclRXpyC0/vHqY
lmofV6/w+aK75rAovllSlfUxrK4ibiCR5IX77hDikd/i0/SeASlBATbUEmK69mZwhFOwuI5/49kg
9Zeb2swW7Lxyt/jTxRcO9mN1qdd0Ajq8EFxgiYwk18qLGXlYF0WvRBR/62MQdUviUXNbP/hcwYLP
KWNDeVjyZk09YwJHQgLX2M5qJX5k2mpGw8igLda0D+HTPcyNYMMGb5IZjMurHc3Z7F+2kbVDOUN0
emrgrMpsQTucnqFuaEDlwmSDZbdjJJ4s76TqT9A7X98VF1Lfi4cKnHgJupI4VTLCoPiIVA7hsVRX
V8leB+9dbogQ3wMBkHzrhyI295yrfZKWtk0jjIiDXIJZa9MtgftOXJMoJdQEYiiJ8wkNbxcQ55TD
seOreIVKEooX3pqBUr5uBsqg0aCa2KRpAGrJJ9Vh597GTorVzexACe4aQm3P1jAT4Eehk513Loix
UFeagNqwd8vGT2pfzqXsVEhvKS/6bBkxVyWEPmR5IbUXi7TTvSPW6ZAxjqPOgejx4D0719L+hKbj
lO53EptGg34r+ABJ9Om+6LLk9al+49LoMIVYHXlOmiYdpnbvQjfN1JwCzr1JOjFNzcJSXBPkOQo3
GIEiBjYNa8g/AuXV0Zo/h7NwLvNZCy7Kq1h8CFGOv3Xup/R+7z+OlL7wk0KdbVMG+8XlLOPVfxQT
YCqMhrLua6YO9cA8noYsVoPIYgzGUTRC+0/gxT4KYjsD4BQFplUe2nXVNeRB8DJnpudQbXGI2QLe
7VAdVXajHlO/LVwHDDvLxeCt/aG6lqnRmQWZLeuaFU9l9+Epg7EjhtMTTEImtULsXhHTz8h3jLet
5XKxnvAiy9fFTvRNu4UbWlHIAtHmlF9C1ajwornYS3enQDAiWSzyjN3a+3MnsDZR4zOkCDd0ORap
89ceVJTOziqFGz8JbH26ouHX/hVTjlpg2d8+4fI1xYF6aLJuDycTUQXEiOwHCTHH6an2hxWgai+0
MWo4zM4HbeIdIkG+kF7sVFt222eukI2ZCt7XmWZmQ1tk7pkO5BwUMkIZ3mMFZr/Q8lFAO3RCSZcj
o8Msx19FuNCaahNA05Yh4e+JzSsvTMBL20azlRR2XNWFB1kEBRYmWpzDNQ4GTF4YZ1kKNv71gZFk
gnF2/ZbqQQ/XuoBVrPDk+OdzHX1ts1gx1qzLWFphI4cQYx8tYPMt8H9cGHzNHHx1TXlAGOfpvnr9
OwFexXX5gx6QocaT6MVPecxsRgKIPuK8r4k9SxLNSAUe0HHQCFnaJye9+QSA2XMraCSQHaVxFumT
UHwGulP1tdOR9hirJ42sqY/fxEjJiNXaj97gveSQE81aKhKJNVyiZOYje+rDiGrac9aFbQ42Ifzx
nD6iRIjvhzjtHh7oCfF8/Mf2gnBu0dfXVkwZ53iKefysrtCtkXAaLCA0jXF8rJZSjAictb6vvR8z
5cgVVvsTe33A9KBHNCCzFv27UXqpxru+P+r0MXq6hQTOoWxxOss1QPn29q2pcwpixhWj3uWgQ6mO
HRt0AarqYdqS/aRqJ/Z74Qk8UfPL61XBbiqiasGiaUIPecOQqUhf91m5Ft3tP8arnMagUxfITLp7
aDLY/MJ0WrejK3Z55IAGnTIWaHl5xUQ66JS640nORRCS4z28bX1O2EKkW6VDGR/c4SiK/y8q1Im1
oNg4hkNyiDYhN8sPXVu2Z66ApVjxq3EYEHS564g25M+vdn+B6AXZYTYM2XN7Ippxpm20NePRClg3
WMUqZ9PrOErklqJJP4lz1aekXojBGw58j5PAJPVXw75aAv0Bv//Wgr4iTK9ZxWZtCPhxxyhFDePy
Mzn3luG3xT+Wi57m7WCxLKKf86YICowhiNLoHWrfBrA48NrGtL0rWJTR6LoA1R5Km+G4uvvU8Es1
blIFdqjzfwprURuH7/GtPMnp6h1+h0quCMD3TCIULfa2ylKDk22klIn1b3Vq6xeTXppiGQwZV5XC
NFGOu3oG1o1nFJ8TF1IjwweABIwuCe4AbeqgzMy8Nj6IYyd5TTFmdvKVnkQE0TjvgIBoc1l5Zly7
O2rHTwQX2KW0gyjzP0EQotcP7kzbQxDnL2JXSYTNO58rsSETDEUviUspKghgQ7Q7biSTr+JYJKmL
zFlXFWBrfh9ERIPbVvxWwnY87A5VWXpbwAM2o/y1aQHYzGZyofwqg7PFUvp9kxlM3UP+pADQGoHf
8jbjeURYqF45//oaSr0J//CI7wEJWaYrApIolCYPpDE+m9up8/6FDYsczYDYkSdisYwlG5iPbBMT
Wjz2vF4F4CdpYaSDNUaU3LZkRrW7R7iwfJzgq6sv7S5pbc61PDyMDQ65M83tUu1iLMVh48cDqese
z9XUq59/YA0gtv6yg5NgNZ4zClY+qGEjVtDwgz0ZVo3ngQNh+vGmZ5vIbZsTc5KkohS1EjlMQw/W
7piwnMqjLB5Fw337T5p3cHqjLWYXi3bd/OQhblYfTGiIdxQE0F41qbX3NCszpXJ/uJtoHA8LGnc6
eHmPZnOFSGndePE6FUgcEf0De+7M9Eywyw/4GbMgC91TzKGn5QGp+Se/hfEITQ0AIvcdgqxOa3IM
pWaVDEQDVSU+bnqFVALClPrT+as2v+m1/kjRMJOu2xAnyjyoPOddo+JCw6Xy8bOpgttlq1T2cwCW
TCEBisIF9lsg5dFwGg1V84H1dqAN0H2ZKIEzIrz9MjEZoJksBKgT+aK4EvlnPk+sAMgaDuvoZTTt
AfGDGoVh0GbHTlVRT6xu00fXXudbyjeKzmOPBLbSlJXilaJ6ZaHbpLAmqLOJ8cym7+zTLShGZpCN
fKSm7Y8Dr1PzEG8Auk9h3ptHevmTkRDLMse56oCsmNTq4YRSyQrXKWkYUiCzu4v/OrL52i7EvIHm
fjJ3Gb2TkVziq6fFfNZJMFyqYVW+4kh6RmfKnQN/V0Dt0RAmZcW9VkLf4t8RqUTIrUsezqZle/Sa
Rt1GRjb9dilZMMoX4pRaqNIWIYe/hCdstxQ+lUxiRShSD2BcfuPOk/fxevBUuDTPBr151Gqn6tBd
/eqbbtvc8CKmApDmqimgwjprXhBLnaMztwC91jLn6khWvsJ1YBZVryMaiTla1f7Eiht2CHZL39KP
pibRkXWN70JYGt0+ohysHBJOCkBbR5r45FwPEvFQE9zJQtAUMuylSKS5hznHU62Ur+l6fOrICjX4
8hVEdoxkUxjNmyZQe3rVA+G7vQ+7sAGS3ayEFH43mHNlq1nTw4cJ4RanJhXjb4W7P9mhl9CQuTlm
2omPq9Uj3b8AnIpUlSOSqkC/lHdcPFsHbRUFALqTZ8iFZdhr7+sL9LexP7eo8NaUmbbkhQvkmF4z
2S8T8LLCCr197ohG7uVNAVfeGBox/TedS+O8hYyaI+zo0448m0c0uhX76cfMfTkr1vmeKc3opJFp
ydw+ixIoCUYhxxw0jv7bWWG2ghAQyJjIIz43L3+8gkIF5HsKZ6S6+kjhMmtTG0ziNZPb7AS+OmOz
xwqvmyg3vNRkRQBrcaIfcpwPaG5TGBI/OdKOFozyEIuRLfepRjIpNpOW9LMvNEdePNwLuBTmP2Py
JE9bQxmYjNtwq9pPYs5S3vSybBTJZUL5OVguwFRu8s2Xw7X4TmuHTH8jbTHptscK9NkTBf0NSkD6
B0PJwMg50P+8ToliKI/1+VXN0uK3maCWX5KLxdQ3i6WxGMeuAIgFcJ5lgLplM/Ob/lwOmNvJiHLW
trgg7ZOmE35BgS6GWm/Y2xLlu4DB6DWAlKI3IVH4mZhfa8RoKEHP04mZ+wILSQNdXL1EHMpwKZZL
81oK32/mymuRp75oK+QxQoM1w0Akh17bZBy+CISsL1ybt+LGaZ0cDdCw396uZFBrgjrn0EgY3JLh
RGh42qz6lO2BthJiD3doC3IkJ3wFL/jvqE8Y8yMi4Fe+3tFJgxMQB3IEGv6Z7Fary++nHaJMMivj
4nZst6u4ezb6hVWIPaMs8dvvqym5NpkuXe/JyFKLQAfZxP6G3owwTL3lgvaiWAdfwnu/B2JysBM1
DRxTJ/5fyIhf43JLImLNZg4ypUTerAYM/RHPsK/cx38DAvBPMyuoPzLTqTk/a/sfCi0GltFrfCAw
8SW82KapqaOgRHM/UPvdRjgWLuF0NcyD7MIzEkId/DGDfR79/IcOc7eqBGofOXdf9MSPHlSLZxR+
Xb3JnMye7ltnjOYPjiMFP71IyaH8upg8VFVq3gspb50v+i8AYnCN0R3H5RQQzB3DvYuzc5bkdwuO
/gK4qwMZoJ5pPaMNrpJBfOZ4BaZXcxBWLtpxeqnFEvOfDKnNXMIJCGfSJYg5WRXbW/HfobsHt2Hm
NJs1LhMv906HnCExUJt91pv6payNuqzUtiHvgo2bcm6zxjXAx1VWcmkKn4wURNjyZdiThnKsQKnq
3erNsc3BopVVhmyGSMmNyazvODTWb71oifs/hUoBvUPzWAEulEAdy2T9c6zupXNBL+m/RVqhhZMr
cmU/OnvmfB37s8c6LA+CB3FNhruvMtwBZeIBb21BovBOuedqk09RHmlLpBep/Sds79RBj1JugWSx
VDCeKj3ue3qWgZjwjEIjOlW78LPadohJla2tJiOWgICwbcdj2UlqjaNcG24elnU7NSJ//eKK3srv
zcueMOyEj0nrg/y0opM7B8St73Q+cYA31HjYMxq1zNeH9vuz+MSgkIHhdnAYaD9aEH7sYGd1scJF
ayXtPyfgjWDYSOWGP2rIl8k4p2Ab8uuMrkaaO0eOBxSgsz5YgbBHINXl+2q9xB/wMWq0nCuo/F62
1rR+PopdgqrbW7Iy5aS7AOU0dOum64ITeOy+gz75IUyPAo31JkMVBvmG0rtmztz3Iq/MVbfUgSst
FwvggAK9Qgk0/IZBcwlQo4n7L4v1261LHm7cJZvob9uPF1k7kPV3XmKUjf92uUhahiSh3fNCEn3s
ZinvV/ubj8sJhDW4kdivA3MXcTaGjB+JMhCgFFE9N2CiKWiRNtIGjsxKwE+FtBHG6eD9zzhkMxjY
mgh5Op2kZ7eVivKF+rmJmFWjRpO9nGrybl4/AFteT86a2Eg4woR0PJRkRGf76XDm0DVZVq/LK+5x
7MQ0+x3TSCvPs355ZKmcq/eYjrMmo4OscPqUAbNZAfIAFvjwLNp8JCd9aH142fAJRN0i4vIk3sHN
2qjyfdo5DLvqDqm70nihBYqe6FgTQjvZWftn77eqH1+1vsKiVkxyGAxJlzMMnSkOUqA9SGVVykKR
x5igAysSfoYZC6GQzeSA9Q8DdbL/E4yc+ijVMtLDQn4FQJufdVpdaCK7sgVF8RcLrbhjz6Pt+lCY
Fc2dPek6wugejQdBBijXd+VOcetbKS0vKJHH4KvlnPby8IHIveOttZ+WBe2NDda9giYtaJozlIbU
8anLyqir3WO7xSYaD3lJMSPRCf2Nq1XJWGIDDzK/mS8KHH5j6tDVRYbx21Ug/DmEtsm2i9zTfQSR
JyG3KzFclroZJp1x4uUF9u7FGWJcyBgiK9s6lYnzeyOHIRsc73C2Zz0cl7S5xcnu2Vjk6hhOJxSc
8ha73r8nI2SB+8Vj/oBHYycPhGMuhq5Bchwzbq5z/YQnYNHR8+gIAZNdaQNcIcOYKaXvaK0B14Xw
gYvB+D/mS+zZ1qHA1rsbH7qaVItr5NxFYeSpNl4lCi5EhI+hh1EaP5QyhZURdOiEbZ4ri3Zkcn0m
hQVpPyyKAtD24TtcUY1C6+9XEleySGTmjuXIe8TqVhfQZi4kCeAZYV6FUIopTAiy/3R3DDtYH8z3
yoHv+KTmA2yU3JuqmXBbexF1rk/cNjsEENUrmBxq3GA7D2nA3PAt6mn9dTAl5a+oZK+u0NOWE6cr
3w4cgzhWB4ZzT7QUKYUwf9lS1y+HXQ/00nVt88MRLvRc91cTdUNE7crGV4p5cVN3Ev5/xeGCv6HU
qTeZUvVfiVNopq24jO5bHUEWBT3Acx14uP6GT53XexVlRaJPPs62cKJX0RZQkqVn1UoWnoVMQGkR
EHZwj8Js9oC/SShy8A2dBXyzmuyF5siZ7JwV406w+BYIyMr6RcTWqpxw4GNDQodV6mKlwuQkSSXO
cgsk+bYEYUlVa1YuC0QGeQ6s19Ubk3xNX8W3Mrg5F6sAaBPimK+88e3JKIh9KklNUq4uXhsXX4Tv
FLpbOIH+PpX4qvJwbl6UFaTw5I5tH5rbQ8PsYPNXCqL7O3emJCuuRCD0HFs2TJVw4lXV5XNqw8dS
Tk1rNb9C4G0ur+fAQQSAE1+foL9gG+2XcQEpsYcaGtaEuWYL7fMfHNIEXS0mZY1h5AOn7cOCzxQt
4D5w+Akemu1fD58fU0BoIzCwACYOMkWaT8UjjgfEOMm7p6pX+CZSQr/LQdf9zttvQU0fmMDt7Nhu
ocnduIB5AIsyZ+OhFmVbbGh8IbAk4KuDLdtUM+eF3dlnjXAL+Hd54mOJxqXKEAzuyNDoRRs+qzsH
JTsaZfwLLN/mrgJVZMknzM+Uyik24OniRTvsrgsmsqymqMHa5ys1l4DpdiAt6y/ii4tYoDz+kdcv
BLQzxHUbWDi60ekI6epD4/fGoSL3Xpm8Jj3Q8Smr9x6T+k9Aa1VEhqXFIcZE1zk1MPwSpEOZTuMy
GwAQZ+1ZBD/Mg1h5OraGdSdWHGxUqz0HD4+BBzKvZLDwhJZbWuGW2aWUYRcMkleK2v3yL9IFsnrB
h1y0oSumNl0ua3sTpoYfY0C37+R131JsQi/DmCF6LTKc4FjFps3gfFe6ms2tESr8KeffDPTAxlkF
G3M1uFSQnFTjAyy2P0cpkif7PgeMbLy6JIE3qoPk58E5qPchN1jHwS5EBFiUbgcb3DcNO/T9T+Jl
b3Vyh/LfOLKK5AihI+lYL8Mu/d4GTScd2fnEzcDsh3c0mzrFRuUshPa5kiAt/Skhrc+P/jtyhAif
TGDFEfmZ+tjtkpUI4YtdSElLiZnJ/fQ+lRSVbhVkx6LpyLr23dWBfOUtxN8h+fY/+AJ/YE/zYypb
nPvOetC7htWRVbtZe9bKfWoZqSjWOGyPlrBKDmcE/HSGLbsCwh9BmSIUZTGqjX4aEsk8hzaNvE5d
zOtzkYkqbEw8ZP+waoJEyWjGC637ifZz1YQZY6xTpUJH96wBjgoHb4mYR9E3imPU3mJWeXOpX4XT
hiWLT9AgoRBjyLxvgNQz4nDoCelmUwsNmaa9ZxEemtgP/Lw2cN6jnB5PdsykIMC+is0p2BU9G+BI
dPBMyMAxZ4qH2MiJ/eTo9nQkKcnH6OKox7KdrRxbK7y9r5Evlh+f4R3OfPd7D0e0mU71WJe/aAD4
LPOCgnJBZ+l2hI8mV45IGjIJNQOoF0JQ6Hx+pL/tB1alW7OBQoOC2Rr89FF1e6jW0Dk5vuEYcI2g
q4XJCKvralCGcQthFyQQTRqucPjg7fNSg2vKaK5CO4frkD/KWz3WBzAJGAh2uFwAwqZFz8IHWy/6
gymTfzyePT72rLpLlG8KyMZeiHF6YZD5st62APEMMiMiOrooUurx418zcWhpv6YGxSAPGU5+V8sa
aNHpFLxwzyE65hyPlzzreMsKEP3hV5u/MVuGU6iCN+YExQTAoVmq5fev+1ZYjqukNhJvqyIfSVas
Olkx+DUveQX5P786STMyyE7GPAp+BsTqb6pEw9nCTrgIhEJlEfnVy94hcz1VJqYhW6jXaZVOAF/L
Eyk8vU1txNYTGJLuZVEX+LDPawdubXWRh+/6a/lQGgbgQizYmh0lLsixprsXS5CoYCtXw3B0LvuJ
8SydTskIQFmzcF2sFfZyNhs1voqyXLnSKJY70/d3QDeLaSIJWS6N5JnwmDk/ny4N79jQKGbdHypA
rByUsJZWf8Yjeh8wyiACalBWR0sfUkg6Jhg3mZO64rv8g9WbOBAYhh+YswmZS5OOSAMjjUs7nb/C
Zm/R7XR8mo/ameCt4d9h0eFa+0A8HQu4s8Gdre/UXdkS+v5lz/nAfCHTNNpboqiuKQP42BGwGQN2
DClqog52QpGVeXrpduo2bzhwz9041vMTDFmnKi6cX3/J2Us6XOnc3bRTBKpGAx6obYU5dIQTmBcY
t5nhOK/oukV+beTNP5ta14H0ibQD0oSFs+9fziML7u0kgDhO8LLhDuCHl0su3zxNMhfJv5XfgKlj
oJXxf3iv7ZUzsXbIIZ19T7Rk/bCqDNpIlXvm5MeNw17ICJS89NWD1guuQZ9u8s1IxTs6uii/tsWg
12o7ZPlIZEsKbb0t2O/5J7jiB7f9U31H+Fep/jlUR0AojRRe9THJVvHhPX3jmtbRjgYeW+/PC5Gp
cGBsFhvcY9vrnOZQNh8oFyREpmuuATWHVGblevVlj26j+5Jfuuv3N0s/2g22rqnpTublsUuto1f1
X1n2uJJWaLfZ/iALMZ8TETWjEk5ZGmtC1S+oUImjcbw5Y4GtgaMAQHXjyvaxFEs+w5Mke1wmthad
j8tZ3OT99pxPqZu0Waiz6G7Y/Kfvv4jVnx+Wo5j0J8nCHbXt20xVjFGdynpoD5AMm1ork0dJI/Gb
jnhRy3LltTzQBU+kiXoVS6WnCLARIdIYHRJJBYelVaU97v4VirO/Hvm3n1r0B4qCFq9hUCIUPliy
y5SHG58mH6w5xG/UiMdAq+A/2wyodp5TDMpfd8BB2Escy3HDe1PtvCUhal6/z3luXNyXoyl7N0L1
2Fw7SPPWpEacWRz8gHfTJea7D+lUX7nRF/J6Mj28R5McuNolQdm7cXBZYIf+QSMrUe23c4lITI3H
fFGjYpBbk9LxBYX0iUqjXCfDf8Pyu4ehFnz9sQSJa40LbeBI6LIUmn8Wx2DQkgB4KrVR+ohRFK03
n28bwx+A222BobOMQjV17dtU9Nq6lI+C/0qTVLBxLTfzL/8tw8IA59TBb/XpSWEY/9dQ8TcXQ38x
8qSfGuwcrjBmGtfbsBlzRuv2BvhZtFlR7Cm8VYy4w7q7gvyJICTqgAsn3T1j/N/uA0bVeFDQoH7D
RSh3XUeyvhXCyCQCboFbfxpl5HYVlhNsRMVK8Cwv7PmTZkB/wRV0LPStn3gbc2xgPAD7mXlLGI1s
fXxoNJov7AsB2Y27kG8sJIdcOYMYAQ4x5IzX3Wvv6Hxh3le3nIXrKVtDMcxIxc1Dg4zFobsdbCmF
s6qf3arzGrfmn1JaGkDxOx251gDeTRr+U3zlEBMDw/o4pOtar6TKSoHuRDcFR0UkQh+qDT6O7dOy
PWtM4T4G9m7K8z/bbZ/BLb9y3/tU65G40FIIOnib3PhBCm+pxUyGNHf1QvJsduX38ItIL59hsC78
Dn2IoAhcnSycppXmqq/9LkwctSFNbrXdabIa801YOPI1/BoSfop+D1219HwpIE5tLEBxu/36x8++
VIjkdynP5yr5zKrGx/DC5V4b71Cxjnx36yBpLTsWHnw8eagl7w1E3egIOg+i9He2XCmLeWoVmG/6
5Pgn53ny+b48Oe8b7Vf6aKEFqVvvc1QJ4rz0czbTe2848As4Ct5QkENqZ+tKFmFJJOKlWLIq57+N
2jN2PnPP/rPr/GQIMRMw4t8662gbC5P7hudgFGxBUTHRIi7uVXbP1fOfpY/7d3EaAv5cMgUv1IYk
lCHs2pLyj99Lk1kZUfvfUHiTgq+zghOuB4/sIN9p47PYe6CD+Gk2JvgV+7mo32W3eIiB2ZOMSrDJ
1WZCmGzcdHg8BhqwfhlpDESUyed+i3BGd6y27uCydQjA+xU/r1YAWLlCaEI4I85tpj7YyASFqSv2
nS++fh36GlMqZR+NWpzu0kBDbJHF1ZhZPBNzKSaqJ8+X+6BqVK+1ddnfGrRgKjHAr5+J4M+fvcP/
042GKu0PMCMF6N51fYxlDoy+Cr6C8duzoAXMGIM6GeIYReMm0qTqApNRZ90nhVojdhOM4SbHTYSo
KniMtFIkajKt3Vogur1S1/u3R6unf1j4dd6cFjYdA49FkTnpjwQfoEk6UcuC+HN/O6Z6CVt1PuWi
RrKzUbLo/SJJg7SSRvF1Y2fuOk0JytNf/dWyh6zjVFXmHL51Qzbcqyl9EYEV8T+6xlNAdyQSUC/4
vnvWgnsHJfhhwROJca1ffzxM6kriGKmSF1OjITddBITg2qkvx8unpGWIV7AiOiIlgyjdO7S4ZqIw
AaY9JcH706eqSrvWg4Np0kGCvNfCD6pEz4IUGUOpbNjkOHfCs8Qj74g4VMuARv+K4f93rK/nFdGU
FeIfd+22c+6YOS+U4EoAP8ZqUhI8FhMc1WHjFQMSHyyVcBAskQ9ZcGucZOfPNQS4QkwCVTh+5f10
wR/aUszfdQVhrD+G/vR2Pd0zZu3yEv8+x5c9n0Nqo5pHIgdMHiUlE76CH8XJGwj8rwUAsGZp4Y0V
hHfMcS9nNOH+fSc4RIFGICzATqjR1pBRPJPTIKLfsmK8R/W402wruKLQXNeQbRagSK+H+USR1PXm
+Qx8ejAT7TLrddDEIGT/MolC+ywo4DRtEDRTqBW84xrRhzRp12PMOvFKPMvsS3Xbargae57WoNyD
aH6EiuqO4NwYcPLwawPLKZH1T8UEa7+851/SrADyUEVK4ku6ZWFq4i8DA4XNunfZY093cm4MnjUj
h8T8ZJkoPSB1bxzq7wd7Yqtzj2VeiPBKIKAxTG+k4tf/epZsVxG7ZX0n35Mvio9GMvxbRYfWWFZS
+G1vOTrx6SHcqM9rPIL5LYh3+nzZNRS7LOQ28Nn4ql5pyhTztwufy6oZCxXQID2CSBA7/5AOiWfh
18G+U8KZqy+x/zZ/jdqjPWgFcRxAvEJXVrf3XLXUzXriL7CXATp0yVjJpLQeN06F4H2PWEh2eg7U
o3RIhV7vUKpsBgwwcfOQcRl7+ztf7Y6z7oCev9TEl5Sj01jbxzA2+FvQGNqeYDESUn+Ig93ShRKE
uZlZv0nCzeKRf6alpQoPqhP5tBRD9QIftQws+AzQ7xKsHMft57b3pR9lBf7DEZObQmPsXHbXlwhW
SdVLv7J5AR3YKYm/KWgO/fufeyrCIz4w5wKt7XlXYawjx0PvVv7v4A4Q1bBDRd2qgrrFSvp5OvS/
UlaDaF3djWPgwLuVu2TXzmAZT+7oVq8GuLfxvy0RQLB1GCJPAXBR58DXtQuBoUZ6GciGbuoSFQT9
iy8NhuGMYSwlJobGiFeLaSkJ6+rqjGI2l5U1mCTc4UfgeS6kyP8UocNQNnJiba38oWC2qB9pY0m1
DyQ4/ZkGsxwWlk+bWR1ppdHjSNSkHBuNglj2W2ERTaFEF7/jSMoroEmxEkQGf9ZmiF3sDLh5XvN/
TF3izz8tfq6m17WrhHhoMQOhZ3my1S4a1UqatIHxvPc2S6L/SV8xv+mF4bc6qvQkPvcHMpiniH6u
GqS/GxP/6ceXfOE2Tx+vorMDgsmVt9zdPlJPd24akCZVcLsmTITcR+b9ZHW+zuJnPWf4LDa6SMMk
yQfkLyLoSs6u8WslryGhi8RnoBZy6ejMqjQ0b2uvpH8gdALwod9ssAbqKKS4pJ1kDfj6rBUrJ/Ml
hA38XlnnfRHUG79qQoZ3Ww6cyBY+KCtZVggUJh1hS99PtZ84aEYSq70PrVd7jKuHHd5HoGax+jEK
uBzj42I8oi0vZMi5psZZsF4C5Ozw3vDDco0kNCbRGq5kI21d/nC7W6j3fiJ3LqRsDcDyrLjZfmNG
zVHxgtgyb4iFgbMPRe6+4ZWghI7x48YukD31pjYlwc8fdxnjb8e7tdQwQez6lX3l3CurbictyWG/
l4hVQ0QASxb24bN+WRSbZ//rCnX0TmxE75HgtqRj5ik61RDG0Cp0owOy7xVCO4cuPXHQr8x7Fp+D
LxnLZqa8189LWv/N6Fe3/mVjafXTXB89CBrZdNH3EelWMNPM0QtsbBEUkNg3Ci8MgRlG6VdFrt+y
px/tcla2+D62MQobK33fOjNh3egPv1NPzKrBHknhP7hvIo7D4cnBQVJnpU8RWmfBvYsF6vTF2kEQ
8Aej8WTIhcllecdLrqmePPW5mB8l8MbteFwd7BaNGys9RfSs0FIImT2RgWR4LwOm7WzwtX/ZowK4
RBr+YOXT4h49TF89nfY4Szxtx4Ex189jrJ15rAv9B5erUXiGKyw3HRKCCis5lqbHgcUZbcIokPQa
KrRPyiVdcvpFdcaBoLDF9MPzLuX0xHLp1Eg2QcTz5DmRRMLaYGlO1IMpRhH1vad8IkCZz47537wY
Q/4gsMR9yfPbmmBW+jMNAOHffT9JLtaoHNdgErH1+ZcjXantZn+I9cZVn2f1p4Tt1dF51mhytLBg
HnHmla7T9x2cWkhUKTcTtEN2RNRMIqrjJMWLEJJJ/bJUHNRqeAeYbm4rZofiAId25JT60ixqNri1
aqmBBGXR8gpBHJgZfXZBTLW7/n9shpsdJFilj73QBHhIwAgFr7Q9y5PaoqnzonjzYA8ojHPgbBtH
CunchSnuWoj27QQDWAB/WcTckhj/oZFgWwyj3yT3tyKmeMialNGXXde8dCJ+Qde0IJ5Z24fFHfCY
1yngJYJTh3kYHstxsxBp5V2A0SVn0fe2TsEAoI/aYnlesFVOL72Vc1XsDF1FNh7/oWnwVJL2/zLC
lKnZlHlx1zfgSO8xE1D7SQTi9xMPJ1+Q/EFQeBu4uMW38QWGqakOOf+J4Y6SYhRny6K0rzt1njZN
Glai+XiafHvQWNLo2Co4lNxZOUbSVPG8qlyVxUzReMTcwFzASzRB+cstUGMKEeNWXoOMJwUQzh0U
JOigG0aW6hV9/+09GXe/IOjeOUl+xSY3SKkrqY1smpZySvbmpTjKCXnrpDBjdXFeV8I54LCpyLLk
PW/ETNTzpIW78jxLABuIzgYBKPdKfeZoQ9YUtundMy3yHce25BBB9PkMMjv0MlFlZwLu57V3Lyef
XLL7OaZv1Yp8IE4+D4Q5bcIeUfMilG00n7hTJveSmlUAhsQOvGixZpQ2zqXeqBlyXlubrAju3PES
nmDKda29+caSCri2bbSvmmJLu9puvhFNff6NfA16MudZmRYDWxsG/hBWnb/v2ZPisus9VgGPelya
siP+pyuqpgOYZc6gQAfcwXKYWlfttWQ5xrIWLBxF7xxN2eRdBjF0DEm5gKwB6zD+Xjvn49HAu+cv
TYM8/VjiJxzVmov5GSMxLc+KAILhQX2hpklKMZC4KsMHTJcqtljoGag8EADbTO7DoMAeUCKFJ3bI
U3sAa3OYmUi5QPf38N9vTM1GondyTkL4AVO7oh+IEFhbQ6Deyme0h6HmSC8EEeQlR3TNhMfL6tvL
aTqFL6gLM75oW/rZ9N5iecDOtcwGHBaGtlai3hxF0yROIQoxeINl5cXOQfkCy8Fbzmhyvx2XRl3L
3vjc43J2jJNCTzG7ZIgkOvpJqfwv0QVH4VDjARH18GFi7Lxa2Sirdpxmi0xPbD5f1ww7jZ8Lbu3r
4Ly86gcOdbfIyaQbXzldZ/XU5XnB+AWmnVgBh77AhbLJeJplTqTQQ51q0KyZ22Bbn4om2CEffXbq
mA2GuSJF7f+h/qenFOXymiVpLNgxJvuX5jVdWlHhkXfdqguLTV9UjBNSt4JCqUc=
`protect end_protected
