-- (C) 2001-2016 Intel Corporation. All rights reserved.
-- This simulation model contains highly confidential and
-- proprietary information of Intel and is being provided
-- in accordance with and subject to the protections of the
-- applicable Intel Program License Subscription Agreement
-- which governs its use and disclosure. Your use of Intel
-- Corporation's design tools, logic functions and other
-- software and tools, and its AMPP partner logic functions,
-- and any output files any of the foregoing (including device
-- programming or simulation files), and any associated
-- documentation or information are expressly subject to the
-- terms and conditions of the Intel Program License Subscription
-- Agreement, Intel MegaCore Function License Agreement, or other
-- applicable license agreement, including, without limitation,
-- that your use is for the sole purpose of simulating designs
-- for use exclusively in logic devices manufactured by Intel and sold
-- by Intel or its authorized distributors. Please refer to the
-- applicable agreement for further details. Intel products and
-- services are protected under numerous U.S. and foreign patents,
-- maskwork rights, copyrights and other intellectual property laws.
-- Intel assumes no responsibility or liability arising out of the
-- application or use of this simulation model.
-- ACDS 16.1
`protect begin_protected
`protect version = 1
`protect encrypt_agent= "Aldec protectip", encrypt_agent_info= "Riviera-PRO 2015.06.92"
`protect key_keyowner= "Aldec", key_keyname= "ALDEC15_001", key_method= "rsa"
`protect encoding= (enctype="base64", line_length= 76, bytes= 256)
`protect key_block
CU+61MySY+d3vwaRARAqzYAlk5MBYpoQHytC2MVTsAes7x2TwB2m+VvVKZlSN2uZjV7xLiBvo7/+
3gLR+g9fvDdT08Pm63suZ9tCrOrIzID0/1O1Ou5bL5L5wXQ9GfEmrBHBx3nM/at+Ob20QI0FQlpz
FytWnnDKungI+uJOLX/hmzmbYYtTvpg02/5meU1VPaawImXPNr+cr0ktP3l84zBGSRqWG9jcXlbE
UIrQdwNBI7QGe54o5InRo357T2h8sTOXXodv2O9vr3wBD/BfG05FTiuHyHPsmTkIO5M9VwwlkSOM
Py06q+W4zj2cdnHUGmVCx6Na81fd6vbSvhxBsA==
`protect data_keyowner= "altera", data_keyname= "altera"
`protect data_method= "aes128-cbc"
`protect encoding= (enctype="base64", line_length= 76, bytes= 114288)
`protect data_block
NUjFo+wysg+GC5ds4VZJ+Kx/BcmY/uqEYUwkYOelsGnSAeBJkfU6MGq+LS+QAGShWk/hJGNXKz9B
osO8Z8V58P0cji0lLk0ayptKSlfX+Lu7Rt7HpPdRPVe15E0MDShPCo6Kzv7eW/yZwcuzWcGLjXDM
JwkfidpAO0JPCFiWOee3Wj6Z/3EwtyE2E030N/S50DU31fZUFUBKo+69g1yI59Hxgv+pFgBZD3mz
yBGROL7CBTunAwFzRH7O6svlJRn4m1LWS0LdsoRPmrf7OWD1W7pLP8yPMbqRIITzcJoPOkvCZZZR
++szNf1xU1eLXWNtwFTl3h+fh4HRs4z6i13xiBQWxSkP2B5OxuiUXat2Mzme2NHCtNTCefrRa7Ug
yO4n9ST4nxbUihtc+K59hm3AgBJeEBQuvsgxmsiDqPuwU73Pv/mY3WLAoPbr5xkxatXnQ+H7Jqgj
jC8xZocLOU8aIzxAytt9uwHeMS6Fgwt4e6nXREhD6Q+I1b35/mbddfD2hg8+jmPiXHBNonFkGZZi
X4HEXVuCu1vKuZ96y5ExyEaN/XZ7LsKs3n71RSjLQFIlJ/ck25O+LkNMXgzKkO9pgA5DgX/Kilib
HZngyLQx1CMi9XplJwBYcaRjeP0/5PmVpziEl/E6Ewalrlqav0jz7M3TRTCeR3B1Q0VGaJ8O5Nrl
+qwkrm48XG8AtVUhHhDHsin7kxCETg2YmlnH/G/WkwH/p9k2MUJQFloniSSW/3U8Sj55FGAhOSSL
TdEg3qTbQ5/fczugYd4XTW7gX9HEDy0r599ZVlXJARyfcnx830BOEOm6tR+2HSXgoadic+QV0S4Z
94GzPysbmq3KW/o4hF26nrrBH0Of2TOkLhmXlby3EPaVkILXu7CIcbSTlgvZqGpOhV6PzsRy0eHR
FZ5gml4Ul9PWm/lmhtSosi/PaUQuxqkrgWAnzAvAT8/0KOIhrU7nlcEaOvVF6QnAm7ucbnKpqfn7
zEncmm+xCReCyU3U3Ep2hteXg+qh0wl7OwfETY2601IU+jkG/kpy5NRltLz2bkDGZxQUu1GnBhqt
MJjRPzNyYdA0f7xmRQBTEXdus0BbgiMEgdLK565/2KNxkIAU53ff3xYiE1TwTYu8SeyEgE9j1rh7
fLp785OlM4f3Sh2/KE++p3nwf06uAOdwp+wj9t3m1rySwGAxdyHmjpNEkmc9XLv5AjS319FB7dRe
0UIHvFU6nLBiFLRjcbdOdPstRYV0SGW9MsvLS/fI2u7cl3pTCIvPMZLaIyWlgOSOb6DrfyFc6R5C
q3A1e0nTs+4vL8yWqTm8raLSE92I6PAMX/wvfOsh/t0lj8ahnLWveUiwrh8Sjv5q4nWiUZAZ3SU0
06DQQh/t5RdfitLRixJ9Si4hn1ZHVvrrzdAHhO+EAXGPxvtPMjFmo+P9DbiW5coM4ftlZ7ag9K5w
B4BOLqIBlQKS1ac4U4f45cit0jqHMbdaxibRCbwy3gnP1exZaMeMZQktEWlCPDYlSc83RHfSJYNA
p3Baw09rnBVXoESnFBG4vI3FfnJBrzDTdih8H++S6dpn5gZpIXsESJlXvwWRNoLbZ0IHF94F6l31
67KZmIb64Rl91jyh4OpTayvUxvwWMMT5jUoYSKnSmvj49KLAlGtzNfTlcXGL76UHLcr5jLbw2oEt
4QRBry0es0LJEN8dW+/Tpn7dEE5AKDTA/1ohGp4ee3KddoFVIcydB2NuC9js65kZfCS5On3dJ+pU
E9NOHssC1W0YFEDNBJnV/3JDQfoTveZ7y8jjFw9UBDXvIyjZ5u+ryVKVatLc/kLXAqcJqim5qrSf
cVJwlvxW5aXBEOQSmEgWDiJ/vLgH0D4OmrwJjvLVS33cvGx5SVaeJ+gqEgRko0dQ0ZA8gNuND24f
BjoPvawu7gfvVouvyHXyr4Y9JRbWvfPrluNMfFv6eof3uOJpL163/0CBY2njKbINF6YGXwTZAyTd
M5bKxQT5LTXwvioU1+A/nenNjN3XumYUy3lzDLTSbwm6M523QdiIB0efJ3UQP8d2LF3Wz5GrIbQT
Gz/O4u94VJsXHlXANnaxoT8m3UtET4ERnb9q3DGtoDz5v8cocP8A1EAogzSGw338Z5QBWHGbHs53
jvX+GjCDTrdqBcr1HX71GfcIRuIIOgu14uDYhYXKrldV3foFBT9aPNlgPWQZYf2+pEDT/LHIgQ86
WUlb5Pm3JPZKviqnIcqpLSpP+OAsnRthfZmjM5FNJFZe49M3glZVSuRIvZGRIIiRa+aYxPEIYOFA
OmcJkv0/ZPf7c8VjAOPLALAC6rhwF+gdGExbupFHR+DrD5uP4tebnb69aRPeCQSgT4zToGmj3xkY
LJmid93nkQIWyx9mzQIlHKb2J1XTu9532h/veGuSNCiGJBeq5NsLMgCUamCHLRgofR9mJq7lnPL3
9t413iocBKyIOUZgcn/0TkONHIIYUkFgUFWo2VcD2oi/FzDab1FtXoybGY22UN1r8tqlaAdUkt34
k7rrpU+T+/5Mw1P8ruVZMB/Oqil+j6fhpgsN6QFe9eAFf33IMtML+1v8TOGFkrcBVRQf5blldXhh
y2LlVWbaJuhsbQOrEbUr5lshiHTNKNblnfq/V5rVgtkvJ2MTJt9CZs1719LKSNYio2NGafoiDDBH
/OEP2u8zuce/JLmlNSE9HIB1FSqo88A0zbN9NjYLEAkabTN9jVOCn772u/wSC2bMAjJkbzX8ASUH
8+0zTFvS4X+70tSWxrtE7xCYc1NISXoawM2LutrRJVOFJtOIqlzff7QHv0qiN/l1j8wi17tRz6aD
8uFwXY+fgoSebJUyyNCxvklxwz7gN/l3FfgoL9psIuDT+wLfTo3o/VAvDhdkFTGG37ovpW0LN34T
YAHrDqrWc2KzXYFYpdBHbsREuSO3ScN3EuTI4rCMdhUKHTofC1FWjSpBwT/bAGmshB5O9/m7gmiT
hzxXmJafnorQAYJ3fpLrDOXJbCP85NE19rOJfUgemk8ZoVoNf+TJT/Joj2V39GpB3J+Azmml02B7
VS9AajOBTpzD3yG6xAOb4u7FPpOz+W6zsNXv9NrQ790S1GIvSQz0k0lOgE7SvHkuN3M7HbIg8aZI
10r+6Shes+IGlrhU4ddpmAnWMUDfMsdBUveRBs1nyTUD1UF8EebvbX9Xhgz6ebj9q9abxtS5Z4Vi
CvpSo/yfb4zxKzEsqOzpjah2sCHIMAOFtnzfyGgxA2NMKHNk39oVBuX/9Sx9qhtH1IHDijay/AAh
V9LSAil+2DSIgixXIi25IcApUWydiP5KOikPxPDCIaIgL0qpoY/DC/11YPR9ENH7IRw3NnuI3R7F
N06I4ietkwmosLLCLleeR8A5ffkE64SS0yp8BlveRi0WlzFNWST+Bf/UDcStTHPTY8IoLRwcZIQ6
fpTh6lspLbkDNyvbBeqYd8Z4SRsfIiGhvrTso+x3xdE7NhTmHpUlyw6nkQVbf03z12m9IKdjixk6
ydf92rnIU22SEZAj3tirqlXGUHd/TNDYJRlMkeParMF3tST4wVY6LxNGceesv6QHH27zoC6GTOhu
hjU3EZyJ11zKSogJCeoyvSgx6tJFThJG9qQgGDHCTg3HqdFetdkVYmTtxRcTMUCUqa1MMPFsiesO
svgrajEkdZ5XZSoI/qXT2T0Qp7MVPr8ldqhWGD4zODiMt1WS8SkPOGRTyuknFUaJK2/VIT2LHwUh
gxzLHnQEoO5XarWq+MtzbJNahhiH9U+3CVRylHLtHuzjzvZTeq9m+sdoa8pXbjuKyiFSgzFdQ4SG
LX7ApJgpdjIT6u97f6P276pqTSdHJFQqQ4y3Qm8b6CNCOX7dnT2QOJWmYHZPHNMplddJcSF2pDtm
pCqNEFIBEc6XKTPnNxuilduds0TBwXuYczqlXffDhQD/YIwYToqxsFbvH6j9bXUxiCoh0HoiTkxA
5gLzJJFcC4vpvXqeNvB8eLFrU7CkhOMrMHd1WSaT3iPQEdFlymAlchvp+lO+VK8BewkvIQQkhZyf
VTYtC1LY/GhUdD5Joz1Ya8yufnVf0opzpopo62YJp1PrnkHHGpCXG26khECXiD3vCiJyMX4zFLH6
csw9TYFqVV407kQQCKke/eGAXvBb8+IrUyvSW9z6Ou1i3YqCWpoLfZo4qa9QIHHRWIIBlxjAyOkd
dmwXVT9Nm+XTNdfAS1OFjtodbUgjvMCKZAxI9eXmNJKfxhxz59MROCD2LCo1capGk5ZIY3sKnfZT
L7OnF7CObaAwejFOCtjh3HdatLG0CSVvWlf/ZP0NfcL2SIv+Yhid10IXf0SWMBt8gpAnZpxV/g2s
o7xcS/qZEmm3Er2jBKvFSZqLC43MSERfiEw8gwvl4dI2IrNkHhHmFFFxVPqbLJBRPvzd6Ab3TrZi
qBIwXH/A4bIUNjckfojNLlqIzF35Desm0d+kzw5y5tnYySBojIXxHY/+hxwsM7C97xGtJXGnIooo
wlHb1c7XGwtNxDBjx1V3K+8ZV+AnKNT5chzZOOZTj6xrx6R/FIfItvkCkq52sIYNiqcSVXwWC4BV
+RRJKjZYTuBU/Adoll8VKA3ynULr0yYyDR7vLLHqVYJnaa4zdtrCNRTx0mL18DlYR/8uEbaVBfsI
YfiTw8vq+VbBNh9K/0zoRxmndRZ3mmsOK7IHDlo6+lGw0o+GP+f+zkOE+8PHtcI1D8Qqri49z+Zs
eNSHpm58awoCYCbeDozQc6tkhIdsrZdItmwRZegORZr3NFzB4X878KCaLWRi0k42S2mwNFLpga5C
w1Swbu7fFLNbbviSwpjFDmAfoLllxLbp9hLH2+fwRF2AOCgLDrBUNPyTYqIjv81wQWa2fo6Btup/
XemSSkBGpCfupUWSZGQME7skdurxaakH6TNP+1KFeNt6I1R2cZGOIKhSh/eiIt1F1Nd7W1GGdvUZ
RK66WRPxXUZyVijiZBUJ3X3qm9Z3c38lWjDis0nX6XAxzioaREgigSjIBuit/Gf6EYjcA1GsTi0E
2Sq0TFEn9JELGoYpNLqinpDHTnUoA8NlIeF4f12fQCV0F3gXBXstcbIR/bV4IYBd+KsEawtMBGl6
/3jM/GE1uatbA5wJzDXirddV4n8LOrl04L//xe6JG4yqXBNv3p9LXVE5JaeECKJeRw+/2sfO3oAj
SLTVyvM8v04SAfE/UbPaL5rNfSyZt2NkE3Z/ceZzbc8hGhqO0k3QgMLEf9YBPG3KcSvhmtGz40bR
Vin8m9ZjPb73P5b7iS2pzrO81eRTokRP9IjiZYhmef5amhT3HXHu0DhJ7z4TtjZNSJ7gXGMmMqm8
NSpdFGMlEOgQA11KY2mKym+04lwmsycOlzxWKGr3FY3NPzXIjTJDKYx5VedNez0pud7TZl/68V3R
Nur3HEPol7brvsJiw3xT8Q/wudpWFFGJU1DQX8nUMOu5DgDt3fX+GlnqqFNkTPAVlBMYclG0i+w8
s5bA2daQbvq16br7uiC14H/N1c/ihwuj3D6BCR+fbCA4AlXRlV8mIB/015kQkOGmQH0S0cGmiKiP
68Wmh/Jym6SxygzpOib/1RMcNNWxx8mw8030qnIeeIN3h6emJjeaYO1hBs4lZUeB8LWLNicetmQc
dXboW1Ak4nxK0Gd74TmrVm/bCHX4cXRfpNodi5u48QlsD3WTP3AZJW9xIICaLDcJ6CNUu/K+YS9U
iRjZKQMtNqRrB5d5F65d1WPrirynFyqfRn/ttpC4zhTFQp/FQXKhNBsK36dvZmJ5AuMlFuHMAksA
YsDJYLj1doRDuhqVqZmfg8vek+57smU3zpZ0A6JOb2sknRxOvqJsGTOPCVe5N+kzvjbk3a1foX3u
1MdrUGqJwypue18Fqq/yFqQre2DtYFAVf70omjrrBF5Tczc7pnAhG14prXgDPcRWK8lZ/C6Vrs7n
OdSFAW2/QVJxZANUCQtNiJWClUjalQXjTgVNmRR367hFcLKdhBgAmfmz08ov9Ud4HImo5nwiWvtk
MuIFtBOjMaJpzLFsv5dyEg62LfZbZmL6/EBZIrQvsHoc+3bkqTF8lutFTjbk6mQc7lBcrvp1tOKA
ddgKEVxFSNJlA87OI5lQcLNqg6lAY3M/n3kBZYn6a1WvKehnblF7IUlCcsYEe0PxWEmp2iwQW4Ky
DjxaYhsVv2OhInRpLDaHI2wPQmvqoFrXN49YAzIVKsE8nVwySvDyLWvdWuY+x+081eD4lBtGPvFH
83hE03DlNjQpOh0txWORDQOQ14ZAr/atBKDBDJ4lFmGrGJXV6GxurUzgqO740KwsYiqo4pM3Kp29
Tew6qjD+WjowcwG8wSLXfyvmfVhxxNvPUoGEzTjEzGpsJCt+XboflrLF+aitfJYAeF2NRB1nEkKN
GtIk0eGO3/dBCuQuS4trIlTKaXhxraU2XzbjXpRbostD78sBzLhNdb91p6j+25JUQN7BO/mnEYUD
PGCVZ75IjSYL+YGi02xm+LRKraaVlXBhf2FuuJUb6st/2qTPZPwvhxpbiDk0RtK+y5rmv8ifbq9k
cIS9C0l5opztBS0E9dr9vsOFkv7jum/gLq9jzqhow5Ka7QEORFP920vuXvEWhJqskw/4pAA9Xmuy
XqAonVhhEwWrzqNB2EMT74vsUQ56l5x/Ne5lcKHweVUfj9DCIjwsLkP8Mxp4CYDsLcIGwiHV5XsC
WJXAr/m5KzWnXLjY8IqDDl0QAfVwMXAtPV826XKBccnEu68B3+BGhRKZ0wuMioPUgL/hffPfad/m
a8hxHrEHLGhgzGI7YzvyHCgI3OmpIocIYzfaKeDZYlPrDF3Owz0rbvjo7V856KZhjrgUwv9mG0RW
wcsRUy+deVKh8nyzRcA4cIGDjrbF/m6bGkCPWSdQhdeZ2yEVfRJazU6+wjTXj6Epwqx4Nfc1U3WH
XUIVXq16rlzqnLSLHjxqId3pDPwsnYwzWewk0YcGI1oqxy46nuOx5FMGbumuqvW1W+uZV9m58LVV
Z7yoxwtPtfwctPltOsa2NKOmjo1oYoqMFLDAwT5lGpuebdI/DDXTPNmsyRrwOSrczT/At489PZn8
SetzWVtybeUaYtNpxoQBtxje/NQwG+9g0YGE1uo8XuvvoBI3koT+8CbHre1bFkaCx/fgoLwse+xZ
Pn0Xw+rSG322S6VUOIL6aNB6Cerotee7/kX5Mi5bfZnr/sJqQLcWQ3OvTPoD4U5on5pJdX91sVfL
qdYkQmhtwRXRpXzSn2nFz9CwawGj0vXyxSGBM0a3T3orhvqcidwrFzonG8Fbc7KYBznCo5ecrPNu
1yRvuYBMqBzDpt4CFEHJL0xhn22gGhjJrCjCH71CG4qIvVh/uBfHJChX5+q+nfEG5PBbxyeIVVCq
dmnBwx0b/KHgu6RmT4bf3E4Dy0r7vLbbJTEFoZO03bo1+/Rizss0oOnD5Xy2KDB+0KGi8GEmUX3M
rhuUCuLac+XOObBuzNwlFH1S9R/oRCzKcJ7FfMc3WU1jJzBgEDHhdXL0z+3zniWbaKgiMyFys14X
Q886f+4ObGXrgDsupipDG8Oq6gURFLndxxJW1wXODiKTmcUP8qolUbt57KgHz93qgURYl07wnH/L
bP9K7fEG6WLNzeKl6LHymG5jsfDsIfmqiteAkEwCiNWK0KbkZZC31hbf+fvNY3D4bQRDseLlyi7g
ZoWd/Drg+e9BX9zg/6WPDx6gOzMaAelIlb74S5FBSMBd2NbCyON7pVcpk6aQuJTjOBfmqUP3hoUO
uR8ooCSuORAVaj0abm1UlZWA1LUsQVSHWInsd4vcI4i1QvHSCp/NNv+ikKM2HvdzCrloFRkyN3uR
E5PSFz32hccL5rZN5/svMplcNjx3+Ywx8Se2wDNe3BT+BcQ/euFs8Tua3osJ8TKzZ+9ELAkyY3CB
Bt05bIvgsU0quEZxZx1Nxmo9cypgvXGkBh8ByvmK4YmtxK0zqJwYD7R9y0SVRtLayHaRNceJDT9j
IhrxyL5klvDXkU3O7/bgmYAmSgL8ECPStqdVFhUa4QBB0KcAHaXCUGAgoyOtfQjC6tkk98if0zPw
KXesyEFw/pR6PdWC9vdDlQTAav/hv8FKlWQZzhXZGL97IDP0Qx6FrBUpi94Dv19R4EVqqQVEL/Ex
MSX95DJrehySeiFXw4Rf3lqzAR+MqQcyiB30X3ujkreU2Lp1H/x/DUBwFFp6liAwTjF0YTdCFPJ7
740gTp8tITiQlQ25a23/YA/GSzpE4v8/2FZTStCX+2rap9HEFj8W4HRiqL4IgovfaTaz2HEvA98e
oXOiPnCqmQsYfDedOvlHhLnxOy3VjtsR29+hAy70oRncYPmTGw6FZEUitmdYdr0CCdDhEky+Ioar
werLoIdtt/TkwQeRcXgYUP9QWC4lOI6l8OONGHlscy5PXAyEEiICHdFKLAy7b3muND1/Fd2ZsG8q
Zz927ibfseEOgbpw+NOUNBhL1mA0Rr3FtjbDByKxO0xvVubfqSKGkJnkCl9T/vHxnMrnPntrImHq
YCGlrj06/NXeA3Z1GCBiHTCZazBz5CEXAPjJQW2bhUG4tLmNNHL5UFl0zLtYv7NXn8Lnu3PyLnK4
r59IwQsExweXvTBrLiSO8wqY0VUCfPAfUaQCNDhb0RtdRrTfIhy7XEgFyhpUm4F5UPS4t2teVyw/
/DA1EuYSi0nL+PeEP34EnMb4xuXT1jgMhWfPWdyxoK4dft9dmbwIjXxKI0yUwOLO8iRURUMwKOIu
U9bnm3jobfEZKWLAGkjdVuZvMsh6OvDtbdJWZWfmNrIvc8vcAwuT0qAcziqDzCVMatS9W7zE3D9B
tE4eikrb3JBZ8IoKoSlis49swJYQnHGgfQraIXAOUq5ExG7LKCJBOFXZ6ACrzgoGSpxxxSuOPgAE
H2840zmPMM0oBJZddpoM7SySsecZ3k680ERelby2spuhHNofO0EWpPz+cWn27fd9fcdsg9S3/Sar
WypwRlij8u+UwsQXi2hN9rYgQa1xObo972PGiYEBnTw8B3/whwCvgeN1DqNNYnXtBn8+ckYhLG8h
SO6CkugoSXJ7CfyO7DkcMXgMsSpXqhAQeYwQHj1FnBhbqKjtuEKqr+ByNUjh9APsOQM3Qz03sPoa
/31f3muCyWbC1W7W3q7IJwOTfKQlJO/l0HAYK6vzEHpNilTLO9G7htRNYoi0nyPypCFs8/dzhzkW
2u1GP2ulJpo1xKv7EfHoGlzCygXvSOyGE8/SREFhj2FOe2YoSO6YManlIRwTQaaDF5EGy/IObE1b
fIgOTjH1yY1/X8QNS4IjaFABMnfUb+XrYfxpHzFp0PIzHa/N9loRysQS9i74Rlxmp8YUp1qlFJby
W55QLOeR9HxPiGsMoqBbS+cODX9xdfdUTtH7OvGAVCEfSlhjpNWSLTyTW4wFY+ucWQ10md+CSn40
aL4b3Rlcrsl/SGuHnFx109b2mqJnmB9NFr618ygFqpDlL8P76BSKQY1LlrGeDI018kcD1Oxn3Tm8
tEsZsOZasVDSt/LbtyMit+kgs2+67fmPtg7BGPG05GZLeOxd/Mfhnfs11ShyEIo4Y53mBIM3YCAb
G9OJcTZ88L5tG8eqYTU4IzvTKf741KDO+i0IMpBJFZBkxZUKeXBdQDo9LOFrC28DHs705pLApNi/
7zp8oTlqYNYbSMwGT9y80UY/O1yJFLJbqLJOVjciWtov/ySHvmIUmIzM5v6ErM9V318pHHCa9jj+
aletxYv8o6fo4a3EqTZzJ4efHV2Tz1fANFomvXW8f2eKGZzznlJYfWPGV1Bavd7E1JvN2PteMuKc
zV4D3DfoQ4Yf/6G6/JEFyqRM0kesHAmF9gkapXv/9rBwjQanPVrwd7Wnd2pzt9HUP8UNLYn+6Iam
GThkYkn8U722FEegaixQyn0E3FzgMf+9QMdWMYaFJmT5Y8+VcZU2/i4mpbg6PjPFHvdUHUflTwVT
16VoQkFzOs5kpiC8yu2/HhqqMfkcNzQsg8IulsYjg3dWu7FxdD/GJnN9Ogk8BSSrinp3Hwnnn3zl
QdcuBsFzOx4wokOz63pQkZ1fbLYbfwEL5Yaimz1TBE/hdvv9GBKZebqCCuvJPR3PdSPzqcdo8a9e
2TlEJuwiQCiLGUu8JBvm3n9+UNK9ocKnrzV5yuAb/DyTPwPSbwZMO5M/bnau9gx6n6cZY5vuxGpi
igYy18Guy/gk51rF3PCUAPDfBeS3EPKyudH8b2Q0yiw3z1KcIe7NlU7fEMyxc6DcnJlvLIWjag8A
5w/Om1eqGLE44i/ZIfWkxq37VI1w0bOFx1ZUrKGgbYjnu/V2HQjiHy229bjf9UFK8ZRpnVHyGZZ/
OY6xyCP0pErznyTjMNf6owkhGrR9pjN6sNYTLyncclT9YJObY5RLc0a+wiuuekaCbqbQkPnvXl/p
kDggt+jHK9m0d653pDsqUKstiBga0in8vOq1ZPuUvoTG9Y7JrAOmlYfrwmsnHCMEeJ2hJkHUMZqa
vnmcl58BgnohdzqmlKHlYrH1gRCjQQ5P1Ggg2ZXfnuDTXd9gRweN7Ig5eW+9+MU8v5VD+SStzMB1
kEvjM1MTq0Reulu8/hmC3qKNE+sDA72jZLRHKdbSaw7uuHECIv1n/dcvzGi0i33xJERN6vwUQMTr
rDsBocdneaNq1G2kCZuDEkLYU87LHzkieAqo26LT9u3iEHDvcLvtsgeBxMp0Dq+0gD0he6fiVc5z
s8DMSdd9RlZqKHgBc4eqew+4IW5SxYHj3Cakdlk8scf4RdVe+N5eaSnkB42xpwdmFdT3GEbkdnQK
e6dilVW5QF2tYmTjvAeuz4TBwvJpkWQMVcrP5/QgoPupkaPzNxSbsticaEOVwN4BJUTS/vm2Fleu
cPaiHvrOch+VJ0BoGrUuToGIpx7wgFqD0phSAIbOS8ynyWIbI0OiN+o9FADpWpmj84qwDkapcMVV
RRQHPL8FPyS8fcHdMkFOUN6N/cgS9wewzqAVorRF1MmhBt9anuaUCT9KSr+gnEWD2Bfdk6h5WqfN
7pdHPQZE9rqBXm5Xc/E49dTCRquaNRcrPh2zywbVeSxt3Hh4oc+SJ8MJnhfNZt/PcBbgebRJDvGR
67A0Or+WPefzs0FQCDZkeu6dWY1gsbKXUlQIf3nHMYYEOunsyq+xA0qqpiWqqVKNat6VhTZRrKNs
KOTqvHhwgz3Qiw8Y2xLC3SqZcgxqBPKTfnb/sn+7BnX+zZj+Q2aWgPyKKH0C1Rn+xQAVaTeKnYm4
VKwAy0a6+pUrpec8WLTA+dbtMb7WLqMbO4NIkqcAHpp/vWRMq1n/EiX4Pi6ItkO13iIXFBtEy0Zz
45w4an3qA1WnjFgvfpFmNaPaRMMotSpNV/rwc6FwGBsscdvmyzzQcn3ya177l/lBuBBR+xO/IMQi
9fMAd3A/7QB4U+4Dmq6TLM+n1r/enFxCe9KlXG7FtJxwNRX+KaJfwSq1Oi87sEPEuU1YD49KxSIH
7V6+lBH9EuJgCEV/mH8s35JJdW+8KG9cOc2ZWPuNy0SukrgcgLYFupC0orrnkYNPLrR3k1o9dmVN
AED2WlIfV6jTVBP72jKqtEXV+v8JaZbE9aVkhQs2P9escuRpu63viHQNFLNVEP2xhYv64EAAQAmb
xjGE1eHDWYTzabtfXVBbyHXxHUCQkA/85puh+vo2dHjxlhFasozsNUjOlBUWb42FD94bHg6PfdF8
AHIGROAyyqaibv8LX6Ej+nHByYfx+9E597IlwIYjjqsQDg+0sX4vdvulUquN85rYnVAD87ECSYR4
VLhosRFF8ZqgepNJ6sYMUhbZy0Wi2Ad5h6DZoUZm3dW+oOkdUmUpRls6cPAbRFul5wB4kWENvLPy
PoFdSwswUZqQEjZ6F6fj2HtpzQuRPxXBEnpNkpK9W4Z/XmSRoXbf/R/eQAjL5h7zI9a2PbP5FgAm
dydkJpn7VD4i3oX2KWOoLdHRsOZiscA3NdAXl6dbp+g0aZtc+TiU5fvMKWfcP98ERFohRnWfr0P/
gSY75QCJi+y49Di6SzZzPMt+oPvpABWzCNCh7rGhEcc8cajGwph9xGuOX0PqYKMTud1p/gdf0Myp
6gh9gYBC5j2Ls2/hz/0WrThI3t357meKySS9I28j0ucykeY7gRRfhnQ/7CHXcinA3uQESz3LV1NB
K9KikWXCBrXVRDrtuNx6a1fguqpqUSUaavIa83kKnGWV6v5XGlEcJv9EUX/7pK6IGUh57ufN+dj7
2/mBchquhOlWqzqP4QKN39jRynKYK8DezMhpJf5b4vjrJAN6DQlUmEGadDQvLX/reoEtoUn6BTRN
EMNoqECChC+cYFh/3X5qokFgLgAhAc3IDmA4wTsLy/fiHXjRHgwWBi/TWjNuinVicOMVmDZqntTB
r/b4omNW8jMmoAxkGQczoJd4LUWIs6mPdf/84zBU2WfkDtm8vmvcJCSOAhRl0flyBD1FpH8zNY4K
aZzYC+JjCvIknX7XLuxMzzRlUpoThCFPJToiIHsCv/0L2sbP1tK0o7AvBWny9fjUfyYFWzDcVe+3
6HR/dDrjOuxSi7Z3Qb6vkheOc55QOacGUXdYLbuM0KNbG7IxSu4nMhufWGUOF6te9XfeyhKQUHnb
/VYaJ1JS6xfsL8nt6aJP3vAIkr/ZDgmSrHnJJnAdXgnwaxOs6KwyyJMvPTGfkW9njblNA60eSECm
f09EbVhCyLKLky4QJFJk6ynExbFDSTzl3+lwfOGcTVncV1HCQ9vP3rvMDUAzbpZTdaR3CBjQ4RFL
mAbMhy/S8ny6iXb9z+FfRn1p3cvs1ocyF2LkCOQ47pq7TVyg4WYwWO0FWPA9A1F69P+KfQIThq0g
gp3EOZ+/piqC21LpUHHwiZljt8GtHLRXf7O0A/p63TLGta1rMuXv1Gqt4LcmuQf43wYDRhVSrq+2
fBOfFTFdhYXy6awIeyLx6YV3IqZXrWVNbN39+I5A1Zob3jUv3EYoVU2GdlNJiNj+aQXQC0roy8yt
b9DF8CPq/5lft1/+S2Z8hRIK9Q8/ghgClzm4xiEh1snnRATXltYzpS3uCTV6QCVZMp8iovhYSKi4
Hh7e5KwVnceiH2Emp2haqROWD4fmNBrM1AYuAtjkUB1xS3ppqNfmpe4WedPoneTi5Qso0hO08mSk
wRaBdXiWPsxLhmD5j03uyKI8Vd/SGxcjfmzfN4XGQHd3EGiG7ILXJFb/YtYm543cCmsyZEhF6wHa
TXMXcIBDO/DgAGmVoNmc6RCNpZytgyGRFIbng6CGGUzFHhAcmxbGxYXp0RbgHggYpsCgOb+EjfC/
WvyGg8xdYSCBHIGEYIrTW7SSv/K8r2BQRqvbRJGblPwXq7+0i8n3uPfifKGtgwf1rguoodFkyo0G
DJ6u6qFDNTO3fuTxfWfL9+hqwZ1G34nh9IklZJqvpzjpERyasSsnQED8myJ1MCOcFTGDrPNNcV9j
/huOe9iTHc7DYpxe8v7f0o0C7AGiEd9MY6IW4R5U5BRSlwmOF+enrrs3TR5w0BBMggy2zFm8WytN
otb7FiicEL4Akp0TAkUu1I0P1RZYKdOFQsX5HLZZFKZkzDEkLEWfJzzRi59Hv7OcOfCGFoo9HGf+
VDcKK2LKJTcukPwrq8PtrXIzrHvkwVAh/w13kW0BdLkYmG0UOnJUzq/giMcHqq4kFXzyGD4Byw8B
1zpyxz6jFUIUSsE4Em/DlHZYyCpqr1ahUKxjZYAzWRYUx//ECQrOJdyASmtiusxywfNu83v6n1Aj
QlrK7D6YK0MUUy4xXsHqlnyB8avRDHnpZ8Z7AZaSq3TjTaLGR5l9eIdu/86FkEpT5SdyVXd3cY4L
ohOFiSQW5syCCQhO8LPFOgPB7iua+9in4ftrcQhnPwK8d1hXtRWbIH1gw1D8smSv7XcJFltVWYv+
MQeBSdjmrFrnEggnBY0LmXe4Mpzg/9ynIUTbvHlXne3K8ERCWD2P8a618fdxVb9vTx40VWrC0bVA
bBMupb8M9WIco2SvtL28JG3JfNVWw2QnrmGz0pywa9u+LsT0aB8Ydj9qtaZNO8Ux/lvTWWmmYvpm
IIEhqveGKEQhKT5rclfCdy4TkxIiprn7eFw7XtK93mQlgQjYfk772/tTzPDsnBKomhQiYUVL94mN
3ERyfVBVhiWE9Y+ItcVGfjOzrPW8s5o7HxFN5kKtUkr+7C4g8iGSYi5LRdrHDnAoaGPOpuDBFiTQ
rdfxIV+P+JkEt5cWD6cbs1mtlSouJXDRHkhz/TUeSepKMK/x1kR7PccGYCQ9EHfNq1yfpE4a1ct8
72z4bVMFaMKoLxBA19gPr5YovDPfA6tdBB2z/Q5qOvmGavSGhYI7Z3sDq5IySTQIZeqwwgv5HW4n
83SwZFUoeX/3aCBoekMOJpKN/f/JzvbxFCxS3m5nGse4EHyY6Vd25EM8nGBoLy0q6m0yKqFLd8z3
/k36t7IkrGXjKy7mPkdm7lsYUX9pt3KAD1JxRMXYufAfXI7y2mg5KmzCJhfXHMpT1Y5PQ70bZ8XT
WYDXH3NZvvPvsHLvljine/78ZVT0wtcYITCBKtdMrJ94glU6xSgviYXgvo03Rxtuwdy9djVrwfKe
6LW2zLxqMOHZEMKmzRTN64eH+jpREIC4s7K3LwwkZVmLSc2HsgVkmUVreZzXnM9q2VX4gLcYviXd
OkAY+hMQMajg5JvpF/xjyTNi5uMxgqrbf1LmEYCV5rz3FSvhK8sS+HzIrOSLd0Kj7LhSdHQjsPXa
RWSHPGzQ8JPI5IsjcWccp9LHGTLayk99Yhw7/KRuQyu5CSJTeWdAAb0uI0OkGyJFh0AVxieIxn95
P+Ea7x9FQ1eATNa4bYPpOpd7owNYsHmD6FqgD84ew8yDts6SG0zlXUFRqQ7ffDpEUOT3gdFzQ8Cs
4t4efUFbevizWT7MMpAgXff5FN27veV0Hz4jWvNvfPnzf3GcGIbF8JkLHn2Q71ER5q61/xcv1HVd
qXaZWJ2EAmPptmTlxLwYIEYue/1tXCtwnZ3pmXWxc91bbESPYfH9lUYvHsbnwWlz1oda5SZquia6
RaaH/6s1ZDB0TVDprTGP3PJCuZk5GfG/cs8hEmUflh4NevKrcKEnW+5hfzfEM0QUkL+mf47lZDX2
9qhRRY3SUUolDh8ZSV+BmV98AX+Oc/4+/73bdCGgxVrUccGsiGC8U8x7bHaBERP5et9hC9Czq4Rw
YDAdSjP4beFGW/VB+WgiMkNh+dJ8oVLE0y5Fg1rs+Eg0bcAWxqQzfoRMCbNJHFjneBNGWwMKwIef
a2S8Jo3QF4+FWm+yNkdADT8x9V/6egpN+UxHhZojmOa6OPb22jQHNX7fT4TCKBDlwLwPyC0V7fam
cFab8LJDk6SQzudcyI3VAsRxpS2hBGcl3SJ1T8DPI064HNeXt7Mk39TIKJNLXzHZ03CbGXu7NgSS
ulBDmlSJsPpTRVMSDfCGwaEzSmDdteaHuCAQqIYafFmvZAbpLGtvhS+3JEoLw8J/Nf7k0mBMDiwk
lapDjCD5MjsvjnjQZ3DmM7qTZy8oBJFZgZIJP0+W/nIqsIiqu82aM5dcXWQ3kNGQPhV6ENH6s4U2
iyxYNMEv5CzV81m/FSCS0/CviWtXPFMXAD2YYoIU6KVZBHVkHOLbctwqUloW7eZpwmKwhvF1Zc31
2QpVJ8I8SLWitFQ8Pg14zIwqdGgr7SNtSRI9kGz3F1KVUH0mbv9cQqzVkxfVI/WODcD37Ha3rNV/
2V4iCAlj3mBmKpT7fnRGDwvFRkN/rZ3aKY50hWAwPRtEue/WNTisZwqicvXPXV7pbrrkLtezNtU/
pKF4fjl1UswSAopq9VtwMAQQhMcxHqgi1AKQFvt/blDPk3rc0pl+N485ziwVdyYwYqZsn08ND8P5
RRDSZAxyzqI0Co49WDMi624CZ7+g5gesqDUC7MTWmWpOTFgL0BKlfY37Nbe6AXAvRkAcjUElpBk3
4hF/IJdN67c02nsPVbpqJ/R87TNb2NuVAYthVJaECjtNnVyzxL4coB+EkmDQQNPdnWXSVr6+fiOI
8XmtruD2MMT5+bcG1BrXe8fq9qqY5P8J2dA34uB6jxKHXyBXH8wPkfDBN0la1/vCgsnrjERhacAZ
rpyJPhPRzYGVQDkg8uiftVP2lH9xMQdYaZgbJLxtDfCC++TzuK3f+MQEkVWlHEXOSy9QJf5/SDj+
q+8uWKrsRLRwghrwF9bRLUbDQ8sg9YUEWLh70g1M775x+7bURm4baSREvK8A1LteZ61w7GTzOjm4
bcyWM/QBGYeq/pQRFfAh7CBFKLAQDeGDBJ0xAKB1cEOZQ1vJh7ye8UocMtk9IwkXzr8LG4MuzyiK
+f9ZEebxp+OFs0apybym+I0uCaefepWkw+J174rchyNV1H/mzu7WdS1sQuNDRNNnHydQS3gATMVZ
D9ZsUclreSCHoSQXEGJketvPwE7zpHFLrkXApTbJ3oGFZyXmhl/nEIdQtYGsUvSlTCDNrLfLv4j6
S6Tas2Eb/+p1aG5z6eGqR8mzVnVS8me6i4k4p6+2C4SZp4GNe814+qFNQa8k2AOB+HUgW5JBy6QA
FdHmyp9Y88Jfn64GwxPumh1Vy4s566An+uokzkJUhVm7/8PGtjCZX5NVZfqTEfcdnPOt0+s+DOBZ
NJbekDbY+DR88eWdPmpy0jo1JyVg0SQHQ5pa/FrC/wctuxFdCEmKwLNxtkx/qKNXLZPcBQ7YU9nU
EjJGSUEC0DBF5u1gZgrJGysob86EAxGa59SyPi/nBhXR5t48Pqb9PzN9GshVNxRCj6Pez2O/TNbh
KfdgUW3hqWHT9u6f3g4Qeaw0nQynT1aZY2FZfDnKDb7E2uam7YUx22OVA/OE0iDcAn05YBRkZHY1
t+XCTpBHS4SrQhiFUlDjQT3iUJNTJZC+Tm+D8fYZQS5CiluCvx6XzQmvKol/6d2Rc6lnO0Em3yun
YDaDnNwBnp/zAyHdEeY+dMLAEPsseIbqfzylQE89n5A/vxGxStcUG1KO70RbEgcLSw1fpBeaL59R
uX6TdL4UBSXMYUr0FIEpYLPK0hGR31KaAlbgSMdCJjgroLIEsxEJdQGRKtJhakFh/d4NqWqaK3B7
V/vTzBD/L9z2k/jZxlFjSWGKN5Regt5qJDxBtgBTLs3BXFnyvXETyeQtbWxLJj9gdE92UlI2Sjsl
LaMZ14nKeb6VsvmG17OEXQ3O6c6RXEKsItcwTOrjQlSusM67RxYtxPRYafu0aV4ObXGSz+NSs2s4
EF2FK2qrnlvkwnnaR/I6uifcHcISx2p1A14c1yfhGktVUSKMswB2fLV6Cp6bnEj13MF2sAgxSVvS
9CQr9CGrdW+sBR5dlGewFUduj7eQesLFlZoNMk3Fpl8OPJ++41NpfNwmMKRdHSK3ZM6ybf3ddwyL
mN5TiTITLqVkuK0izyYQQKz+jV5LKtt5jOH+BQogEupZEgXkBgMpZos/fj+6j3ZrdeUSVGCoZa6d
8p1VDSMERjbE3Rvc9I9naTJyYRhULIB+7hyP5p/Xgh43KJKv1jdXMwtoUxM46iB2PD4wMzc2qZem
ABqVJpRogINnb4VFPUDYEpoHsJpr0dPialV9pNxR+4CUXg967chiFCnHPpgaU0JvQjhKPf5ZRsuy
nhrKfA2RWENAjMApaUu+5G4mkEv9egeKRa2SSNRloDEfofyDh6NajUMyrDqWvA1jK8Bh2PVrFxgI
RvRzOl6z6gIfKRe4lOSqXWW+uH61Dzfh5H+kh1qCrh3pT2R7DhLxCO3X8qAsCDNKToa8GP1JRcUK
8FpNYs8jUecOkpHLekHnI1tcAiyV9Arb51McJbyScmnC/ZsdOhFFHuJZNimiUJ2mqa7YQacsI5/Y
/5nGvjXe+J6kfiQSD8Phjzf8QJPARZwLBfiRC6gI7tCStVuUDweWfvJMo+r1sKgpxZvajGqZTOyW
5H6MaC+FiApjwElZtsCa1R9d4rwGnezmhfQijR9EAB9SR8tx/E5huYsixqV95NaTI+Kk6dzualzi
+kFwF1yPbhANjeZ4luVdo9rwmpnJBNruVoxqcG4161fXOw4cgsJlujT/mK8bvV6qkZCSgg0r2Nwc
1ll6TErWiGueFAZr7ScH6vL8SL0vIztg30KVDvkCf0Ms4Kdw+Wttj1p335boG7qWaGw1WCNMOwIU
M4aCFiIPnOQ66HO576moEhGbZ7dLUJOTNjrm2RFoFYB9zh2Z+wfHOh6BhnSwqiADqZjTyokPdVM/
BFjCmajS3MUxBp8jO9k29BUShqprA6AOmQnuImH9VvWebOdfVjRbqV/BlV+ohzhG3WLWFqayypw7
hiH1jJ9jT9fQeBqWsM7cuPmVZsx1MwP7iab8epzfhwn9p5i+euh7xcK2r5H0aSgVL0fkF2ZOhDFl
fP3Dk+L8jgpLPfgQgstgBkW9AxmPUxOWaCsFy9yBZAoNEGcDA0+Ok5q1d2r5nbnVEeju4XYK8TQv
M4EgI/yAQ/zL7bxeomWLhO/9AJw9AxQA4QY08h5J6p6zLBYpEezYScmpG3pMQEK1v1V1zQFakNOc
biUiZJYO7fy6JEN0rGig3gAblNQjB8vLFeMu2U1YpW+kW7tVNU6C0uR7f3OGx8D0ucGj+d2HxPVN
D7LTyrjs/w2KGmaYC2qRJPCMsw5OyAFFw1en0VjJPqxkXWTfUxKRE6ib5oC5VJUwKA7YkjOgRddA
6nieFnJAk0UpvJYoPsam9Bv01vyGD9qlGnMnxmo0QH2qEThYKxf4kHb8FC3XXYZ6GoruUhqTmwY1
MaO68vns1l46aBovkBMfIJLG4OdOL2lhDKHtII6evwnjGvaFj5WtA3HY+fU14feUzIx6+3JtMivL
8COOgkrYM5ulxj9QIJe5VXVALIjpwq+oja3fAtkSfU3ZA0IJc6n6yVvilSTrK2q+qvl7a3mtXNzZ
/gc3hOZvo3JDUv/bRitbbxTUYjPBL3Mqr7FJeu9PgIAR2UoZEqfZe/zEmWXNs0ljBAvfZM2mn1lV
DaOL7RqkcV0mBMnkZvdCBM6OBxO4wj4ld2XG4p4tSlorEE7pEFbh3kcN29CFxP7SIPoBl50wX44k
enI+Z7W5cv84m3rJ6WEtv15zptNMBA+oifb0iSROPkX/21lJ0ySxKhzQN94k2IAwzUx7SCmtPGMN
0b6G1GJgegpgwiYR+r2UP58HSBufzZ7k7luoRQ8nGeK3MGPyre4wLxmOhQC8wCdMrCz/qJ80HXZE
uvBzeDiYS9ILUyB3KrzJzwKQncpTccAZz2jRTEF4jcGnVJ6R1RM2S1jZMVNU2kWyqjmCYEW+uiFC
HPa4NalJvfYcjpBxtf2eimBRocpKK/Yr7/JlhlDDBiMeWL2wGMHDhjBikcfYUIe+llRWcTNGOb2H
IM5zJ01PxFOBLwhuL5ggFv7rCt1RvffW/VxxGk4gYdkINHX/LQL0O1RgRB20ux2+l/dGsVkpoTUS
P+CFbrAyMkw5w5scLBBGWzA6sr13aJT4qWuzXh+h2ZmGHRLAtkF/A1GDX8ZOvi6qZn+k5CJbTNvr
YQtAL7mTudPsoqahbnc7Qu0dMLdZJpl/AgQ9gjVKsG9v/ZJ+MCbXvfpbOtGqt071xbOgcjMhNDJC
9DukXKfdB9I7aIRDQ3S059UR2sAmXozp/lb5BpxRXvnJ5nU8LalTF7g7UySXEe4y5mGeMGkFHr/t
GMrWztZEW0RCq7vIGmyq3i1p7CjbqB3zZs6G6BM5jHnha9FucfmWq4RdNUji+/5e033e2Qu/om+W
9LAyK8twIV7TqZg0Ud8epW+QLF93jTa1fTN81eJ+RR5FP1000Bjj4PE95SpqycVlbddYvmw0OeJB
lnl3auIGsCGOyYh2WPNCEIlzuo4fjCLwsc5Z0Qd60NOjgJHhMOyUagIjquQS0fRYKN59P18UQmxw
lSDE2l6oDV7U83HB6tvAT5mepPk8HnfAUDSO/oBvUU3L3aGbiVxJ5yIdNjuq9fckHBtc+tHVtqND
Da/1H/U/ce4zK5DJ+Oy54Z/RN2TkpzIoHLM9iqfDPpu2Kgm0ujfg5HouDQ3yC1zNFu5899ZfifXA
+5884WTF1PF7Jw1PJBQfjqE0ozJ9Y47Jv0K0rj9l9hBwaFx/PtJe2OjCTwNQxaKV+oxqlt+ZSbu1
plJjIDLktSgfDJE9JrrKZD0fAladoiX++cNsjpeuqA9XEerA27cprvhK/j8cSTiDOZJoCYtJymGD
G7vsxLUwo7BDOMpLQo/vovujFHFBaMqsEtvTO1rU9SOxKyTyad/wNZsiW5CPxr7jdEGTbgbqyv04
15Q86AO+RWW3SQl+jAIPVdAlZ0TxYoU6G9FFnLWQ/WgKALBMnMKv/pHECzjOSp/vYzttYkEzSbMj
bB+DWcUVeP4eAMbD1pS/iRlBGSVGKr3K41rBSmFT+JOBnNOKIIxYNMQXPh9Cm1qD1Nzo40W5oi09
SjHQbEgMFVEpo2jpZmC3mQU6NxMx1zwM5jghdr3NHY1cqkMBQzw7iCy4yRuOkDZXGxrTkaX13ney
oPEriSlZlU7GejZgS5HR5cIFabILYgjJFzjVcgeeW0IVfJzWw3p9bq5dNnh9SgrQcElQTpvS1/Og
Gr0d75WCARWC9dnwfT4dmMMAVL4bOOWiBzeMLnpKZMj94iDauIZZFHHP4J22T2SK2+1jFGlVGa1S
sm8Xl+KikEiS5yr9o6G2eH5V736kVA2SENbMtJBR8KT8OU+MNp9DPGFXLeh6s5lCjrVkM2mMD2aA
8nr5QhXRl7ku4MSxHBYEXanjKo5FX8rTDNlgeP/jzLS10eIV+GAlxXMyyk5zJyaVyF20gSdFohv3
sj9HYQq05769kwu5X+Hypgt1iSXiVlnSdAxHk1lz3TbKmBVFr3XZJWelmElG6ukUc758P18z51X4
xnkAFLuvVibN7bOFXnFE3FKhGgcbWeBkPOlUnRkkEv/jCL2bKm8FTQWfXRUSw3jTPq7VXd61g1F3
+/nEPbTaqmtpK5nFgoe/bGCc+zPjbQtuTTdrgTPSBHgCFT5MqkPKbs+JjdJcCS2gRTJR/dZblZw/
NCe3TSAk2xsA14npww6f1eRNrC8tDBv/my0VUQLcjAL6Y6NdLtvVYGVFMXaeSynz1VOuabYNP/CJ
YFidt/HwWUR2XmYXHvx+ppysXTCuaMtL5jOTH/LyRVAuEW5EjLd95mFdBD94sNBqXJHpKCCudqtV
Zx9zOcYiycsu143B4BrktOIoj1eSFrMilFgEMxcQuKkiU8Vj/XndRj4mHbs/RVKo+DIMQ9TL0c1Q
Qb8FxXpW70an5IrW9VTH+DUiOxIc/68DzxKepjSjjwzQcdDSo50x+ZBJdxLRy5ZsxWfA1RTIszOk
DbN/ITcEORbYmVsTIMZXzj9FGQa9Dlyxcx3QbcPlG5niTwrCpYEnCORiJiQX99HSgp9l97HoXGmv
nIP0ZuZfMiZqSCAPb7lOkISd7+sIxbBJOpxSJh3q8+yoqn+Pppml3hVFxA9IgW+WcYT926ANP2Gd
bpR9s2YyXALTh2s+uWsVTp5ZAo3+dzO7K2WPhHSc6pRGeZEImBqRemgP+D+/b1VNWhf4rTk8QH+h
x+aJQRZTH/53la0vAfP2S4oM7Gp4WD/pGWlZbQYQQQ460QA1+nglkNqxx1a54LMKuIDNu2Lf65n8
3hlgk3M9gbs2OzWvYvf5SKhlcAcWNnnnO7BPUfUPAk9unVRb+wfnLLC99GXCrx4ZfxT/M8HuYZVe
Ni15TmgcINlFgan/W1lbQVv8EsldYzVtho7wJGSRndc4S81yWCJ8gwvovWV6QwdJ9HRG15mhCZSG
P6ICua+3awX+4cCI+cUvD2f2Ee1BK1nSLv3iVGaX5lVb3AWL5CgSWnWpjPc3WxjzDovf0Z+KKLs+
rkHp6ZQdW86MMtjlpVsWLQq9QlSK3c0MSLoBmygJn2Vot1t3hJFhB0SihRwAoUsgv8sn2SqB5lgU
2akxvXQCWo0//H9JgC37iksBIvpwqKna1NUNIOVmcr5sUFS2VwslwiMYeJBYVC9IzbnX6X6xExsc
wCTz3rny4m+9nIkuaMc7m0ErZ9KkCs9FzjvH1Kqbj7J5HtkyFb6rFmZ+Dhd7WVj0l2ttcRk2OsYh
4veO/bbLqmuSUV5Hoi6DsfgzGOJX9Yzuklu/avhrbWewaGY68vbHV1nYuERT/jqJ0u/WBZVjydzE
KbDZuOfnuHdWoCXDjZcY38S/N1M95sLlgZCKMkByIBW7NfLXQxXBvfeqg5pUnur2kpk8gcjCX3kI
DleiyfgIRXkyfTXScoHlZ5LBtr51jTD7aNkg4Ebya78NP0lM8stTisUnWLtSasn4yO+wN0EEytTy
zQcFWCmUI3hOFZ7BmK5ZkwzrjYWxDbOPGlzX5guSyLEa1gcbsdXvPTSkVfMqz5EvhMKj/K4h27fU
2VJd6k9DCYxyvFURemrpJPvzgd49QAlThHUgrXS6t7MmGl9CiZ0/vMZArrPpDYZBjvWyXrcIKMVO
YvE8iTP9Z03lziRunJTxmWh7an/prwOs0ApXFWBpm7ls3BfZaNu7yvmx56hFEfPtuIlActlygH37
S61i+ipGNE5ciuZFupKMRlwFDaKFEDawNOFNw/g0sg3DJ7XgaZ3IAxp/MWD8xM1IvXKWjMeCzWVm
mL3q9dkajerjh4ih6Uia7CtzXMMLAoErlOenzcru5nk6YJC1Dh36hdgnrz0YeJuA07ruXwhZF/RO
hVsLAGX5rg5DFdO+Tg7Cwo8M0+yv2GAbR6Gou0kpyyzBq2svgB0P3x1uGOlkGFcNsJJg2zIzUrLN
GAZquy7ro+3hzZxmxTpIS7jkhZpV00JkNqCYrGpy80ZLMVVyWsZZ5kjwyMsUDdHFXHxCHsHe4iPr
wzlp+3ym9RZi5eayyn6/+YEArl/NiBNLNknHxLjdlREs72apVKc+kza0BeJHGGIDjciOBpni6zNq
UoSGB0GzJxbrxRzaB3ct8AScC8tS67skqCIXI5L6ITKQd8GXDu5E4T9VbJqVD0mkxzrn3HSzunCL
iikMzc0KfdpHdBryKuvTqnOYbgfgo7SCnnf8GsjFzVlSd12oOYC28eExQINpwK1h9uGfyPnkybnO
XzbZkf3xLgn+Q1zhwDJXZVgEG5Nt1u2Ul1+Ti3cs3i+o3BcPxuHr+NJw8k98hYeLXmLnz1KspWNV
mK0fmX2jobi4dzr18bD92np6t1teh9XTSw3QjQqA/C7Lth+B8PG9mtTNXN8rLWGYcqRDIU+jRiNY
KLilqau9a6EYC+w589icKOgZo1abVSCmG7+HF/W2xYHQuS6sCQY5/Lev6HUxct/EMZtju/oKkVAy
3MkWhcfhxMI/Bs0FjSYLD8k4qxMy5ZZahhnoiZK240t4nv/lBVbVcL/nWilIq7nQBldnm93mn+MS
NdzhcG4PlEkNliQcfd7tufRXZnM1PiKQtatJuBSp2i17JJPGmgURVjiHR04TOzv4nYrLLA6EYuhi
gPMj3a/G4mSXQY+mr6K5VqXjNOQfXMn/m/x1FPeEvoaxRveT4AuTFkepEvDhVPFQGe924FyZ9rX7
ROgZ6/TQQddfhN2SBJVwUGtXynXSs+S4ak5uwCREp1GCh2vc29IAj9MG7FWhAcvH4fyUrp37572t
IOyowQ8F0PfCzKZYu8P+t8xnu63gRSLlTLidCTWY37y/uiyDGMuQJKqSEC8+2YnA7hrGM9giadtn
m1uAV0QHDOAlWiDBmrxREusEGbPTMGt4VYOYW9TLR/fYIxK2piFrEclA5X3j3G0Fbxy7IVygCpoi
mR1UUrUQ1wd0M6KyKFlfvWyK8nzPX4BKRpqi+PTncNIxoDWYKeRB+Oycp91Wpw2LrTKMGgRaIK+s
fU1ikSelqV+PYgHv4jFUtg6M4sTRm6pJprl6DLuHIe4n2/vWHnfMBdcMwuY/y7SJ4OlHlWlBKP1v
L57DzraemaSQpAA3qkJtgSQTtgmISqXGehzty4qAA2wWtei3cvxzb7hR0Xo0q8S08BZZwA6WCgs7
0IqY2ZJbY32lNeHnOVi9xIsbfjWiEPcwHet/trB7MYZydtMBnFRFTy6KHnm0rnn33od4a892yQ1T
0W3PV6O7QDG6vSAGXkJ5CBNhzc2oFXq+R6etPjU3HUkMcNflCxMluZgGBQn9itvcUkzrLMwt3lTI
WC2M498x4ljEpP1DxNC9/qCzGO9+z2fs6S3oEMhM2pNnraE+7SXAHg2mtGb6jXziUt1H5ixKtRt5
DUecf+rdcQilI83gl9f7AugEsnAe0YFUXXwrqeie/Eb+ofyCKVB/87qwOQ4XUNS7Z4/7kTa3CmQf
Pzx6CmxT6TY9y0hG/VEOvXLjZuhTKTZ9h26/fn83bkyoUOCQIPA3MwnqF4WEQbSDx0ykM/gdMI1/
0zOeM/BUdiKREzIM0kZaIEmTvWC6n5fHD34OHlMZ5w11ib+P6q/xJ7IZdYpfYWf6phssO/x/+fPp
PSyMsFujt2RbfjWqe09yXM8Wv5u0Z4jpGkC5QI5E8djwyk2H2y2naAYsA+is5xcIi3jcpC8NXGYy
r6LBIBHrB5wMOIPvvhpe/xIwCmUR+zMZQ9sldJ7B53D53QEKFQqciuB89jytkGCezZDIf2FIweca
PNnQGPE10sB30DFeaXaAuycSkg6W2bo0r/hVZtYHxN+D27t0Lq4sFcw977uM605CoOlWRdRJU+bn
cArsXRpGEea8zoVH9VuYhhDu2gveQyOEnppDhf59t9gQa2rPBpbrJz9L2yLIqpGB0R5a0BolZefx
xIFSxl4Uk5n28EIDYFOBS7Mfs+F1yog45fjWIdqiYEgfIFsWT8UvrahMIWxcEBoCjsR53VuIBxQw
apg5rBg2ikGIaP4+Z3R0czKvGN8R1a8YLawECXEJm1e99CVOySKH2CLUgBtgt8CnTwA+rArIXzZ2
jyi3UUe4Rs/zyH6PvrnCCkZA9LkrXm2QKUwpEtlkneplDvScWEizYZV6ZmB0fY8MQd+CmOaBdH/n
tovnFK0J81p6f4JUbrw7WhHPhNOFjve4tRZqi3JfJXzjfTyXGPbCjO65Haq/K9lH8ppK5p6LENPY
tvzbfk0It8QVFsY2qwJ4qLMaaijw4RwbjWbbBSfiULhtTjK88kQItrscPIj7VplQTVSdfLcD4I4m
/CW4fTUukkZ1Ec7+UOvZlDPlo6CVwSFUPziHyFyjHvc45FmLRRVVbqD+cVGu15xqh7GhZ8O7q1SM
10/qboIJLiW9m4MpyUBDPBlsP97UjfKPEnCQQrRCcls+Iui/orqif2col1hBZaXe59TVBdNcHtYP
7kgzxYRLWJreap/dwqdAcyfyag97FJdFVxqqYxVnBnhz+1XVrZtZgXP9f5N4wMZayyyTJL97vngV
s+hqRl5Jr9+A9uinzy0S9c5EcaJogXSZAVXvusM3mGyZ50kGAgAVA6UQSOkVivh9KXaWvX82ULl0
ma4QLc5WR8oCK5BfYKyA7l8S9cfHSEtZxWpNdYUfjjzthdNMLAk0ZuG+xoeqrE3wzHbKYvFX/9so
Li9zCsG382rwgS4yBSocxGw58yLvPHV6X0HlXVOVXTC2J7NWGUkULwq/Jg7jDK4YgZywZ2trIaqC
Z0l1024zlIjBT5ld3sQdwTj8LfUk7pYZNC5kqBYlTrgaKbQwqIo2AtxNu0EYfrRi+CfAS4XzxCFO
aH3bEfu/LyPN59t9mLbE4CWeyjITLdz12Hv2irGi0vFuMncTD2N7dJXXhRVCvkZziYwyMzAQXsWI
eRzJSnRhLYTAD7ywclOl8s0uBvBd7Mb4cKReCl3UnwbTTuqYMdnDpEtnI1GSUW1arntXXQf4q+/v
0WyS4h4lz9SxK7P2PGixf5n1m6oVNYIx5h1m1AOppXDO2C58qqao4S9IUDOKhiqTYi7GL6nhZrvj
CnacI5fwcsfH2VSgu2+DG+AdV0ezpgSD+n/eJCOV+CoqWvfpR+RjDYTcrNDK3p9KkAsEKpmOaRs2
4cbyiHqh4b8q5BezG50dq6hz6vWzCIxdiCwFNA/tzAlTDhh5dPdJ+znDT4ccFSU2k3QzYzmL+FSs
T8u+AmWQzzG/iHIcnK5I5Lxb+14Ui1yv5u8i35v4RPIWvGXuYvXrbErdSMu/9uRN0ghovgAyetjV
bubKWjQE+CMRCp6on3TB2ezcTh/anV1Y47FWGGbtQyTizvQqtY4X5F67X4B5ff6lMwmPdyuLSFOm
c6d1sKbDpXPoHkTJ6woihdM1BUa80yXNYS2Y8UwNamYPPrhZTdSJgyiKt4I0zVfwjOQR274Iewoh
zfqFrvHprrVhYvFNnTJCcLb7wzlRI6PzVGDe5zTkduSe981hNHbyJ5N81UKtRtYsM8i90ZzZ0XXI
wRCpL3Ktxtf1Td5TMiusDQDragY2DTAzLM+1yaB6O3f6sO5d1lWvEqnT8+f62H2oAwsG5991x4ac
L50dlI6x4f9Bbl9zTQC4SwI2lJtLg0Q7QVe8HJyoS0TIrC43qZwT+Pj4e+WkXWn5xHw4toWhWSmR
dcNkDxOdnQI9F5TYYMjenzdB8Tinx3ObNtFh+iGSyhBmgtyrXEO3TW7mu5HGvht/9mdJD8cfFgzc
pKxfueYtY8t8IOEKqNMaucK+uAXI4kzqS0viHdSCVlqTPiAwwEJohnBkBHh0leuPT2XhGInV2RyJ
9F6jTfICc3kjUYgFqsKB+1RSgWAxVyj7bTdocAtii5PU4G3r2+1ON/ZV27DjmJd7rYaCVeSAMVg2
yrGixyivVO0WVwTIM3sA6U8pwzaaGhRbMRF5vzFyxZWCjUSSGp/wOS4t1w2W786JHAwH1VQDR7kM
nWOgeLvBZMHrnQFV/tv3LRW8+Sv8bprPeZEd4Gzn8lq9OxPF6YSApZcp/pk2g+0VTJuJTfZiDVdS
guuBJoePwXU0ojRVBm179tWJKHmltsHxy9z70ZPCB/d8nRSI//LaWzzXnbL5KJykSoldj5AFUZwV
AR2CFFzIQIlOiHqZFNGpNnMsExeWV19G+IDRdugD1LFlY8tO5tKN3oaGdZrIIT+ojpphMoKkTK3Z
yGLA92WH9zQsKlmxFCgRU5UGLa86EXAuOSMWE4w5/IY8IKct2RqmpQkw9Z9CSM+XfUo1tMYuENv4
Zcb8a1cCmf00vf1o5EvsfUEAdhi0qU1BLH0BEmahBYQj4k9iE29injLay4MOymjM4DAMBCgGZ/sN
IyjCSUr6l5H8QVtOYnv+QuuZrFK2tKZblyAGmb9u6E3OsRQo9gFrHAoZswWGDAzpY3XqrVXQNGqQ
LPjUAPkBVqfHyXNajo1IriQeZ1FTA1m+tIBslRlT/9C3ER7ojUsr7DuZfge8Kp5lEI86UJAXKR3g
cC0FaNquECcqiXDtPzgjYHztjS03SuORZRJSRBnyVX6jvV+ZrVxXNyyA+E7YmNQgb4GKnNWeJkRz
CNPEYIvYQibBMIEqu4emhhfp8TbO2C86T44WR7ZDpWMBhLb+cIHXpMdMAuhB6qbhVtlBvNqdJ4WK
FaNlX0r1a3JjrHMSBz+4LrXshojlMKhU7amr8X4mwmu+se8B7K8UVFSNklAKlJyZxQ+N2Tryj6MQ
nTlo1sfp287q9VwHfQNpYwegxYAoe7IgcUrPhDYnoEc1Y83+inzULVAPGBc/dk2QY0MeM5Z2z8eU
E+bC8SkhrsDUGADWLXpkTmlbNgq68ScfqwHRfweVFFGefHKXiUEvJDgsACHStAYNSbeUG6j2AOfe
ajtwYf90ZtH1aRIT4JWd57MT73a19oJUspG6Ykfy4gpQTMjicZ5faiy/nHgJm44QtxfsTfT89kxp
7qooPda01JlPBubb56ge+fWeufaOz7YVSYZJk64NdanncjqG0crHL0Xo63MlNtPPFLYiFU3vLuQj
dN/Va9ix5ioF15HCWXpQt1J83pmpLDVuuDhWqdxT+WInEeq1VPn+z810UWgiqgLzzEuNttt8CuRP
FQ5ErWUdfQEwlR3CUNvMPgAny5oct9G+YKGubmMIlW3bc3gGhd86waS6Fc5bMYQaD97UKbD9muGm
brExWYPZVBIcQm0XIV0NfvQcFgZ9zZN4MlYxO41r8D0eJzx2hW0Ne1u7N4WlsOyQrtrr9DxyR5ml
/MBpSC/+u3zWKOs1e4VYwQsbSnERzVQP1Myq1vHH6tR+jQLXNzt1duH+ENIW0utlZR6cn/hljA0e
gBIsZDeYtI4dATkk6VYfb7ObtEH/2++P5ap6/broQHX1BU2gTohCx0gLnXl5FrLcWAypjcJHcqPC
0yNZH+eivTzas8LLPNg9jKELM83QNDQXkttkzi+hoGHzl8CoHIgoAGYioFkoE4LaK53dyq1Kzo9G
+zjUcRI+Nqnq8M9tBaM9CxRTEJc5l/m2MB+GAoWQq6vnpzEpTMQ+GQaUdqNlDeIAVaPO3pA4Wtie
rvd//MYdJ1On6dDeGTNLecqwpc9YkTLt6ajVVL3ye02JgCQj2nwdUQyU3BwMx/5Rspb09mC68q3m
GVamkpbGCGcEJRKfT6arA8azn//3BOr/W9gVJUIouqg52YNMNd95lOyKmKDzGk/ZnWPDoYtITqEp
B1gM0MjgeBaxB6Nqsqe/nCTfLewpVcfNOqneq9V+NXMZBu/nCJ5FpJ3zJ33+DLppTb+Zl6iPHpz/
v4eQM5RM3DVhgy4y2u6XwLDEjBGrW7F4BrnvDKq3DPwZDvBNBQHmvDdAmLNMQ210cWYfTXymmYY6
3M8DN+ktR5+OZdkUs99IWb+YHuI+GZ2i2/IJC/KxZWawZoEcPqHyADvNbJvVV6fSArf3imC/bskz
VCHJanOiHr81h7JAQRr87FLlyW+2U0gSuohGAPbjQ+DZcIulUtnojzrs3tzYHGb9YDqVGKtdtQ3c
i2CrI1Du35B/VITaZoIVPN0dMXDpl1my/+srDdig2Y1Cz6xH3XV3ScCUAR9ohuV8OtFjCyjU37cp
R5g8SX6Xj+dxMoYCe/M+ffrFJ3kUH4czZKrPx4lCNofdClXnusZ6/mqDUL8Vh6oyzJP+I0TwwZ4Y
NoYlTCfPwSgvnGUXIA63YEumfUeGPA4xlAFKKcuIZumnHALITJbQZE/U9YYVvAjyTAidm0ivLz6x
r3fIurv4VExnitkvSrAElV9Rvp3SIdSreO3vzWoNN70CrQLPVsdW9Nr0EEgbzDVYwHJcN4vX4TMh
+/zGIxnnXz5sr1oyXmBwBdf/Rb5VrphtwCdnKnIJo56BPjMCClr52Zi2G3FNZ0BTCe11WjB44KGb
IR05lCjxbSehwe13zDIw/1ElQOco5sX6JmpWlW4oGuJCic/4nBTqPfFFUpRqqyqORaN4LSWr8Zcj
jJDN0BHP9LrC7bhPx9+9eMpMb9VWX1HEnWMJp9Ksi4G2ZRKLWbRpr/WoKJpWrrP8SEkdk0C0wp5Y
7f3jqgDEJxNPPKDv+knl/5FC2gokAt/QBY4uQrSna7y1jABKIOETrhVB9q9NF159EZMEyoOacfuv
AKjvgrp96KDFyYzoQZNtPsm40Tr/8dEIjCKkWR1flM31gbYSaKx02ZME9AzDQqMzLK7z0//r/zya
WvMQyStjzulCyypXr2Xmwb/QZ5BOZHQEuTdsJqAqdLlb9HGyfQUVrlhsaUxZYrx/7aASGi8tIJ3S
oOU8RBi2QKClj75gvkbyvFUO0cpR6f7Y8PNNlpvkYjiNBZ2QCi3jePlfMnh51sKOJHWfi7prFtMg
kBAKRFBgUB+7xgfSfHO387ElC1iXD9HP3HNHBt95q4i2MQsigkv+ZUv7QLMtQDNzBo5NImahQCeA
voCEjMIDszwg9RU8ovH0LAPNIz2b2PXWWX4yII3hGkIrnpwStQZIoITEd693rfizZXUGfRmJ3tRA
zK3deBsZPYBfabl2mpW/gKdVBcZ5vMUzUCDi9pKGOieNTEAcgziICJi8J0EYY0jr8lHD/tOW07RP
ObZ1jQERuDReVB2JEm8U7UIj65irGkYmpC9npxFwxJpwUKf5zLn+yV8uMmltYwhE7biGlTq0Ca7d
3rLCcsWbJejokr1d8CkPI9usd2ywJGoPCNeJAza/d0zahgHomseVrwl10yenuKI67AWB+m0hP1UF
oF87Qxlml/hprh52NF/4IDdhlEf/l/aBjgO3csxGowALTBtC/X6iPuQUiXvEZ9UHOZ886hiCauC1
8lgPNEJWR30+ecB84CI0iX50zAKaiLq5UEs7WxwHovjYkMtJ1knrtCZ163GKlcWxMLam5Sw3BThf
lOBdYLths2qZ8JFHr4nCXMCVK5m6kgF4XTPyZ75T0IxGCaLvkMy8g6PnJvP9SLWWl2sXeOVqEtTh
iQlVFK0s8CyBJsVumaB0lQ9nWKHoPVr8vNfJAB8gbUQx/HC2Plqr34wAQnkI21ooLlds63tmji9A
7OCafyi7v3CG+pr616+lqZ9ehAr3RVwlingM+TW5n6yZln9V51MQRtjChZchn0UQpLn/mC68CHmE
AB7ZYjgdnmJBWl0DA2f7yNgGb5Ck3mBqc4ggAyvTOaJ+fImRPdCJa1In+1/j6RGv2BddUrjCvghc
zzXB6mpIQdMzw+IA5wkEHmZdK5G7Fg1wp0c30Zs+c3BS5GxA/JlVp2cTja+aoC3EOl7h7xVHtJZu
psYQPdcvKPWVEyUmtvZ84OmqUvGH9I0WQFHWsY7tVZingmyqG+wMC5Tr2QnWWWhP+JPCpToPiccI
nerib2goHDnDMuWctVSxhl9jTgeU2fHG1Ix683kxbt10VipT/udvduhhP7YlO+DXbkaXFM1rnISH
TfpC4OxgVZVyu4ww85vXBKGeBMwXFuUinLizLOg/QMNNPgFSt1z+tmGJ7wGMbyEX9jJTcqFNevPA
1SW87/tPLl9Zo3iJRf2jgdsSzAHglmDW9NEvFAmivUOnxek6/YK0QIi/Z+OOj0B/r2EVxF7sT0A2
UtEaEB+uCW+NI6CdrQKlEZk9sapzaMxYs9QH3pISZGc3/qBLMbt9AmhfkXD+irolQjMPi4/4Ml1p
naPl8Rzq9W04GdKz/2eBqe1EhF5sYNmjzAyRCXaSr5F9zDpSrqyLYlgj3k9PTrK067Ewzqi2hGHR
HD57Vf2z35yle+wBdY6RhCd0n3A46k+FzAwJURKeXzGor+1xQlkksOlpNWv7S/DVApmYWbOo+Kqo
uIzM8F57TlM9pXKN4QEZvG+uyDWuaamvOxaRoGOq6oKfp+xIMxecq5yFtf0Nw2nPWexXVF1q2Jdp
ZsASEqlVjG4U19yU3lTLqBJbce7yJDSztYEp+GXMpA54QdiK5XeMkQDBkl0pFcpicV1YTc3Fxt0F
O/jrT1FedVwpdbR+nhrrEvKxGN/nCsNtruaxUJ5CfEb5iKacPphdPcOuOIGpWO8cLK0qTW/Nf5dk
HpHPXbhSDqofFGTNMEVkKRku5DFY1oiZhD3dqS86OWGj/5PnhEAIUTuhCgToVrVEFh8ao8m+RyP5
YaAWtPvHLPUR/vxALbGA+TnEDU7C2OMZsQZGPdiil9+i3gRMJPahUDOaKn+wJYrquisgqo4bQtQi
rOM6zop7TKm7AtTYi34+0Nlj8y5zVT0dcpzlczuuDHp/2abuhsw7K2oNPELRtsn3IEqK9r1LrAe7
FZ9JLyC+xkfdFFdX50WIoRIJCNkaXoC6zQ0tZsFfMJIod0dDhQZWtONkyYjfogxsPDKI/Fb5G5Rj
nU/xGYOK0c5vWBi8+pxJf/w3XXUhUqjwJK3oOyiaUUb73dU5c048aOgOMB7+5I+YWWIiliQq1d2K
TUPh2g0nlQ+IgpkPdbNadLd+on/dokNeY4qpBngFwlMM4cELmltoGRX1DvntoXnBzhIEWUkR+v40
iI4CKcnBtM3sSWVpLDk7qGbO48gyH9Wx4YKCA//DIoSh5TVZ/QIYCFcoRELfryqIquq0d79YbbpR
18ivvNi/ZaAEq9BVkTo7ndjyCOO8AVcbGtRX5ddNZysLqnNliV8f56tuScABDNO6STB8ZPBYKhKt
3NVHjyoTDLek2t4jkdg/KKONOsOTJKHewI4DIQpZ7D6FQmySzRmmrjdKswx6DqGQjZbZFHY9kncN
+ZwVq5M6S8G8h1P/jT1aU3Xv8BPleb5W8R5aW8ApoAFsAUuBEl+zYknFfAI/liGXvYjpi3ZGee/a
fRYodSRkKpmwOZRFxQZZKvSszopUCx3zM1mQ0JaTR9XC6rHTqnqdg06doJO3YolTVBx/x4wUuLjo
u/TX90WnNZ9l+/pJNcmQn+wNpZtLh4aTG2Cau5YaRMeEGj96kZvsImnjP9p2A4+uKjoffATWoDe/
+ieiWkuS7FG4+bn2SpPYTOGZ88S1EZs+iSr8SCcsjRWYV58NkBjm0C6h9Pzfa92aKbMW0qSyLZA0
4Bxhwy6z4inffqZvjPZcr81qABmGixKqccbv2/SjziRA5zhzG7TaKCxdQ/3XUxTUif+6gvb4h1Tw
dci85NH68KLwtcgwHe5sE6WxAt6x6gSYpk3TMoklOkBo2CTgqooKDM0qHHIh1ZagsAvIcQBoLbbS
PKvS485zg8N1fiVTnG3pxMiCtyU2QM8nLuPB6sbzgoLj8VacB2IcYejIHEthxghYBmm4Y9Uzi+tr
l+v4mtGrqa5E8o8RGnZU3rcAZx9oUm1hgTWKts4got/bFI6JunmJhSKUHYX1AuTC7bYGxNF3MKlq
Ry90SnA04H1GHIa2HUqkLLmY96iMAJlyqT0l/wb0LKhyX43E2pbNQ9A2czjGvcsFI/fqX28umWxW
bBbeha/s40udTgAi5TkDkallDgqVej5HcsBAByK/aVNj/FDscn/gp/F8FVaROdvIxIDRJOWB9RTC
zJcSPL6mlSncUszPFHhkZsKFT7B5bs6rvH+0nxU3HvKF3ryoFXiskjbt/KvlrWVgI0+P8yTrZVEv
hOzk9gj+OKY1QcdL2CpPSTUDo2RqSCgdgbfW7lgm5f8bFnNfLN7poEDLks1as0olmOurnQL65R9h
0Dfy4ESDXhS60WvKx2gYZjS3CJp0sAlhBsYo40vLlpeIobQrmFv9MzDRrllsom+Ya9HZf5kP6O3m
3jQa5k2GLj2dl5MQK6Wfxup8yE3uBv8rf/PopHbW+mXdZYp9d9VRbLNSUoNV1DyOV75h5qasrVyK
W8tV7O19x6JQk3wO3jEaq5Z8WumWETjvEy/URhnRk+Dknufg42Wpa4vmaVz2JQgLaQ/OTTYJLKIc
YDBvZrNU1yl1d6/Nozsz+i4l7jQEfuOfEWbbG7qPVv6K7jzZS2cv9QOV18GyULvz+vJ9+cdpc1bI
Cjhox+AFaOesO9e7GPIw4G5kxxjDMTpW/iL5d7iqbHMTZRMBLrpIyoWQcfILfh7/rkYj3lERnJWT
yOLqBy1AgsGnUFlbOgd3HQ5Vjy0YiG9bEvtvzWNQl29+u1lI3R8GZk5F5dNrUUW1EXdUfMxuRo44
eG9nT8d4blhAibSnuVZ6jL7VLww2xJLVZbi3ZX92RvCNE45cXDJbRwjjjHmS9jWV0+UhpUcsrBR/
jPhz4znzj4JdW0a+ZuBu6q8uQWIh6LN/Lf5cJj6zkRKBA3a22+N0XzVIpVzgk1W+se89oI5pg5ea
Sp60h/2lyqylDbKcZAeRtNV5mKzyaAVcDoOqJppmBAv6tWgFvzwhwSyu59QlEPUxmU+mmqWZ7UZS
TEI5fNAIz7bx6rrfgfTo0tjFzTbSKjXgNh+9UWrk+J5RwaUfXy0ru9dFTTRv6p5NbCBScMyhYGl/
04Ccod0wIg15yj933VI0AzjeWZVEb0avG3jdgFkZHfci6l0PRt+0eHxmRWw20cSrLOgrUVwTw3+P
qiWhtIWxGT4LEdBDhTbt6Rq0saDAz+Tlc4EB55do656TvpQHSNd/rIGEb+ZdYLTYBd82/kVFe7u+
86+/bKt820twb3OFmB0phxHT03OhSRUxJh1Hw/G55ms2DEGEuNVgKx+3eAPjZFSDmLJNbEY1N1tj
IPASz0cnZSRBjaRnThS23/gC9KvGj/tr1bmcebsui5WKawqZPgHnvwlIdWIi9V+GFo8pgGHvwuBM
2fIZoFCRXLINueo4TG7LxV6CfJWa4yHSP92POTeUKeeYku3oFhnUjknxIn/8SqCZc8XbAXRdCuJC
0FwL+xMzRGrPRvXkf2iQxluWkWeWQtipsctBtAUkmQy6O5T++1H0y1rL4N01QBw7G3y2FYFWxBNk
BlRQkUqE9LihNuOAaa8TT6uL2P6UmySRiwskDyoBJbnCkUdo0HTUxvhu7IGr2p+45/WE+/fzGXYc
+DOyoArZoN+w38WEVBlWk1uhbWSjlL51ZSW5pgNfBkKPUAggDU87miFrurJXQgKT48Bg/UXI90T/
C6PBmkXGdb75sNDCKczJJPARtdHPPEIp1hQRbWTx17qD0ctwLJpGIoulnkna878lP9mFt/QCftzb
n6ixEljTdA1KweZF9cLWb8bEpawDOu1Ys3JnxtXFA5GrVuPxORxSSzwQxaTZIr4r6UPCn6eEtf/E
+d7lyMaj5wwftiVBBXBKvjlSZL3P/VJZb1j/3aRafAh5Im7PL3v9deUUW9MU3qzd/1RVqtZsBEh9
Ljja+FxIHjooIjCKXR0bPTOERcHr+p4jdg/tZDIu/1gT3IgGhKeSUSgXeLAsKprx7zF1y8jzaPio
M4q0jjwssNmHmw7bKFuGi6GGmRcxNDP0DqIMUQJfROgsuKWE5TTVLApJxAxN9LqR8JlEr4MrH2zf
u1Tj2iIiEacIVlmfxRJnsyM0MReUn1KA2mCoZenFxMVGLwl3ii8pMb2wnol9t+eMqjZn7+kXK3Xk
5gU/rzrociVKUlv2rJ304rR9MF6CvfHgOt5JphNQAwxkK6hMUQs0ppw/rXKiFfU4Nhep6f6skkaD
UL+1DM5XNpz8N0mk3hXMi+gYnrI+Y0GYvOYEbK0VsXkMLr7UfW+UfDKzHFGEY0T7chyTWisM43U8
2G2feig51CIwXuVhDizDt90o84vo0R44nA7yl5lRtpKMtxSxi5mksGzN4i6bx/DOcDjhhLBINnXS
4wk+OjVPa7STU5Rx7CkbQFuN3kjrVi5DZE0Ef/z7mBxdeC9isGK5wIq15h/4SL0Bhm0QFvukISYA
1qwInEB6Loe+j1YG1QWwonUo5ewyB8WYOPXKGQKzcYh+G4VO/iKs6SB2QgnxOnJgcy8rYM14rTPI
3ipsR1D+PQdQfkitiZJ9wptajkYE7/0YpqmUIku76PNxxf+s4j/1xJvIlEbtDhnvcQNFASk2Oybi
CJWnK9kNPT99Bf3FFjLQaUD04+cvi7Izf9sbiIL6pApHF8zu8FKfxuuIQmwa2AalRd/+DEzZU9nn
3FpW/Fd4dAlzWO/lv8leIBuRCCvvgeu6C5G1JD44Lo66dbMZ/K/uEiDQPxfKhGdjivjPx+DvKY7U
7R5zuuRTYVFShi1PkL689gYBCfJUzoDQ4E8ytU28ZHnnt3ZB6ntd0Hnv2tcqoQhuo7s3OMtknzHG
SpPKacanfA9Rz3XsWKfCkMZbzQlHR6XxmtyC4rlNn8ephXQcmbokfCFo0Gp24fGlMSkv2ShfEvqz
Oi6ulJ6tdInnNveWfnK6dFeH7A3OJdYaxyeEdB3rYpc+SCMruz+jSGN7FGETTEMDCMxuQqY+qLSx
dykfaIOzbZQu56jD0fiVjkMjsN9+hhWxwslvxefHHK7LKxPDQ/53tBEg5RS6bjZDheYyEZfCTzM0
PwSLeyZ9rtWASN+QI/pCZ9T/7/wUEh+AtTbFdOlfiZEkuyMiJbRniiDtcpc8Ks0HZbW87Ktxc2i2
o4f1vRpLjNqn1OHicVi3h2IpKKTsN2NcBFdHGZ/Pg+E6TD52VJ0yoOsC6Ed4dcX6hdyHB59lfxHr
4JSYA/3YZExN+F2thl5zcOUvMcPPOR/TRGzBubI6/anV0GfG2TutkQWwptoZ1huXE7zOJrB/nMY0
QeVuBmN9Jl6CozsI8kEAEliTvWis3yGnjc6Uxl1v/G707AWF0Qjgr6EWGPMIkMITdBamoGOebgGX
onrQtcbsV5t1/Ba1DwBXWlelcSSOc4ec+DmQLgDAtKfzoabZhZZhum0lNRGpS+jyxT7v4AHgo+ug
7K1vRUgz06VkoJUDkYeG1nh2g/ELoEe1WNAKSqtZ9Kac3K+E0MBWsLjli7CUNVM4qkMBT2uaddso
yivsNuYUHI3cwS/L/deXHXkSExrErFa9df0jz86ILQp00mxdd90UwUDJuXtuN4nAs54Cli+dXFtT
YP0rFvf7XfOGl3YG32m2NmcZei/gF6E3CwRSikiAqvCYetO2YLUY3wFbIB053RsbGVVuZJmvz59w
7tpxLVC7q+C1L1Ta8t5a2Xbbw4Nj79aReGl4imU2P/FIUmnipcR+zidAn1aXGrgm9KBnldiTMLti
Pasl3S+Z48ADCLt1jzqT5qU42mc6gjXMRwjENWqBUga89ajTExfY8SlwmWLPvPhETlaIasj1bef7
RH+kxEYJLIK9xqqztCFt/VizAz5pTA0/HNRKUkACyigGADDtNNA1SbhbZiz6Rh7U+1iTN5kz44nZ
WvluOHu60WtIIYuxNifziKRdjrM6W4Uh+phJsa4Rm5wERDmLgG3L/nL2K/mVAc+/sJ/ew8M5qUfV
DXNnmDP5nWmV4R+Tq/I7fodqzK5izT7S+OPr4CdFAjPmjeSQNG8zP+nMRIJdgN5pGmDLQ/zXNgvu
vcp8yJ+GZOwJyR8B/pTGtZV4m84JQEg7X1eZIqQpTjpsX1fbGuqWUR6diiuaPhELIfU1YazW0a/0
dJ7UQ8RdlCjfjuMgCbJTa/XCuGMsudCWWBfI9od/UjWDLj6jdpE6dGnHu3e1vEYkvWzdI4AhAykl
B6EoNwEzwS74wNYL8EswfoGjiEp3p4Ma76tVoALzWxw0q1ixQrS69lNXowP4ZXGM5Yg6wADW/NLj
/JUw8BGHTHYFCx8ZsYz8ZUdu89Vgbih+YTbDB6JVo4Rk/3GKvkzlkRsgfgPv9FCPKsZ+zbBiCqmN
2yjmXabkLho/NzbQc0TGY6SxUZv55M5aahoZw+Zi946iZ3sd/bPKlu1hb2v3CEr/a3q6u2vigMmr
JJRUUQ2kLlizsFvH+btjUXZ0yAB2GpJ0HMEuKgq/eh5C0bBmr+6/Nbn4BqL/y639ifgX7Zw3ZOag
VViIEsQIf/wS0QuhaxfDCmchgFQpcD8lWQlVmU6PoB8y98GwqZi1wcHJYYXxWSsznpWyC2FLFGaO
SitD4UUHXSjsOPzUz1X3Pp7ubPjATnDXq/wNyb7sCPOACS1ppNYGzSnfGKlfPvjsTa2jmBulLdli
7hS5QZVAugy7uRhBPKzVNXK3V4VFTwEMh0ridtH7Z/dZywfCyJ0Gc3ASc/ysXSejfmb/z5z1XBqv
VTnVdHXpTfEC5gieUVlTOEzRMXA8ctN5ljqYprR7surfmNLkoKJBGjHVueEFIQDX8/6zpWmxcYRZ
JlufBo0E6cvUa7abyrxLbGLsqDzdTfVSLBC7h5Ekw6A0q9U+42g1NiXHeqIZ2YHJpOGhj3fJn28F
Ihat3gx09xkQgjUHqvhfuxwE+DzSWPEySH07YbPgpJEIbDorHp6OxTuzrCduq6PSFn3opT5OScHF
ygmPu7iw2liR0MlE2h/AMeg6SgeqxmZEyPfvlWrCKYW+Jh9PKBopucr7bPG/NZtdJXllYq6eKsm8
i+kErK97SzY4hr18ZgRRZqXL1ucgeY+Na/WYOzcxAiszm7xmY9XOzMxRe4sNBg1oP8uPEO7ZT7UY
habftXJfQNicnq2xrBTYPzJ1P1cDIi09zqSiMrt9SARJNu4EbYf9Q16WSgKH2HBDL9vX0uQChJj2
P4zvn+Wgg/mNPK6D1zoOtL7Sb/UTFdPKWca9xjhnbmcQKmDpPLgXbUbaMCF0OTDytZBcsfYdWgJ7
EqvNNM97tnZQ7PvWjetIJMRCrbhsg3fwRW957dxtUdv1sECbzAk74mPYUIcQcSKrY/yabmdsFkUj
r0bs3sPZKclloeTqLqoPT72Ro/ufL8dLpQpNJ/b+fpiUzqg9qRbTf1mQQY/tFnTXMt1bvuRepPXP
tpDufj8SvD/iv2kkfCJyNskxN7Iq+VKw582XqoMX1MHI2mnHD3NyESbgPRDW0x60fhBtUD82ampy
wgrRFAmvl869qPUyqz4kBokkzyfNo1tSCiwlB0MjCVBWC5rqyaF50IoEOKRlZ2OIHEHrCp9fgPyd
ZaAro5THBBtXakN+yFfpyofmfLBxRTYyo8f6HtVDGiv/S1hJj4XAcLvM1IBhUxMIyvnuAvJJBs3A
AhcUUBHK21cd8Pi3jkHPPGFkJoUgDa5RwxOtixnfMbfGnFGj8UYEmu1b6+0mNWnvSh9n/dORXi24
716msLBXRwZOUteyTVo1c3qHcLiVeU5ZCav2KJCl+frS9tVtTf++E5QdrGf5UeqIY+CzWf7MGQQ8
qR6nJly4di6/ts6Yjn3ox61TjiawxPUk/LWAyO7rhoVrPH8Pnqvhuh0GRhB9b1qc8agtH8UbhH7k
47CyoCRuYG5YFTNaEuKZXs4/VQmJOhg2pMvUjijf6uKfwBPaARKUBQoW7QY8YytR2ngfxMixqNkc
Pifi6kkn7Q9kLO4OI1f5VBD+zvEussf0mvNEcM2uevRXIJkYZMGkSgeavhPjSVnWT9Bgfi/sswBj
dRTGBn8gUcVOHLZczJ4CGIbusKf9sF+oSgp6RKd8HqDOIAlNvCuaX/7F1BdUZWlNVgey48WNuZfb
7zNCNsPkYhqJteM2HnXCVWCvrnhCV4KWD6s6KGH41M1e41FnowZKtXqN+7x5sOHMJPDdg+v6bFKN
+/ebEl6gqe5PDa9Qr9WJqD6r3/2SVQaNvM1oqwSazPA7RYHhPuW6Te+K3ht91I1j6dw624pQV67f
bZYMQZmD2QgHD4RHNu5m+2zWaCoqKOVik+S0eTVr23cqJ8TK5HmRDqNuOq4kiZEx9Kvmb1Ns6JLY
rbRWBgxvNCWckrRp1EdMM9WKu2jxregOtiUq/j6s9jpF/PVsgfPseQL94vBkFjJqkJHdUjyFk3ML
tgE0urN/3RXjzBokZYv4v2KrqaA8VbTRN2qnCpd9CdS5qmCGAPG5az6Kxy/JWDVDcaMoqf7UpVfA
zRw1vxRdSgx73P2Ca6Vjy7EYKrPc2ai0y3J7EokY2Ydp9nWM00xj2ynqT8LtUWzqMvd2naKDwdJp
Zx2tS2Gdz2lYd9cjIRPcpmOmKavd4cRbr4WWOF/eW+wXjy3wQmpMlztivcJIA/XTzgK0BrYdMznl
5PZAUQQaa9PJBR9EcC4Vt+irk2Jz0JVxVb4SoLE8Y1lKpphYltoJOA5OyuoI16gWA6/DUj3/1xvH
I49mA6s5oJKoZsNAU7iORQfvMo5EVIQlTzbH4sYCZZqTmBn2RQyd88urqgzpYmKVr4FVSpKrfo/M
ExGDI8TUEqV38NoGa7iVsOZzYTIqwnYqh72h+AGs1mEJP4M9BFAN+H1TBFmjYVVnX2wWqgxTxw/i
Pp3MFZugnTJdW9ZhR6yWkdmNdyBbQeUg0/Z+c0kfjgNJZrCA7biBpN8BCd6wQqh/MEO5hCcCRQ95
tDZ4kPY5Lbd2mtgL5+cPMvJP4GG0nuOG1Ic8mbOAKZaJdufT/NbRvnB0wEUu1vo3vyWRA63duU7g
h7zdoh941gT0yFEvjPLwIwJ31f7aIrBSiFNJVQ7qA69KiemzUP9SP1luOpAYS6/xG3q+Mr45mM09
RPFW40xHh5TEXeDflFHSDTmGowM2r3cGLAKEfuZYA1eGHvbndBspFBvZ1GJf8MRRxb1pao4zd2hO
5oKn1aSgzqfVidBLs4LInv+FdIiwtOHv3M/8d9XB7jte/WebQwWDizTN4jxCJWyFUyEj6H+EOsd/
VIovTDjkaMvwevI7Hm1BshpBbfgfY47ueKlLwqsZbl+tRXHLipyuQTuagiXl0Wr9oouUOqcYz7qc
5w4JHPzX2gFA82AMVFFcC2c6FEEtIniuytKJO7ipPz8uThnxqa5b0Fy9LiF+FeCVhC+Sfy2dMXCH
eAiSiS5DAV2ZTndeuzYbwFhfwj7VYlvnxX3LzxjqLElUE4QWaVuGYRmAcuZpsc8NJSS41zbA4npW
BdhW3FxBZ8WRSSuD2ckdyVoimuEhT+58+RWn0U7AdeEEl2eNUIMN+PsW3mlbBn7cuZcYjQXcoOcq
kcSonV0VyB4kIZwPzFDccYh2VqWcHXdBgyhmL9lv9DOCEFRQNIa81ij5daebkFsJe5ukx7XAv5Eg
X+lEikCF7+cXOFmxFWsYpAT9Xhy9rMOhozebnhjyEQK+ixZ1ygmFOxpKROU/CoxgL+FBUlw1mfno
Mk/mdfZGAWmme75dAaHU0eNqQxbI486J7EaLpvUVp75iynozF7s2NO7taHj8vDM7k7tyIwruGNqx
ZAwvzrad5QdQZEieot85eH3NmmFAW9WDzcPs+eyA00fStEUSUloJ1j/Hvhv7lcwvb7/K63qy8lyY
mnGR7A58/UBOgQ1Jk/ONejBfcHMBIp2kA/wGpn1sv/qVnJbov2dBK6sKmubjuwxgJGJ0b7bZBEof
h8kbKVODUt8OpAxy96jQDyI6HiQE7fIHjNkMbwsK2PyO5/TMpovjb9PXdV5zyg0l+jtL/43Au+V+
mbvlbyuyxRjYWiBVXXvuhXqut2zAzFCz7/rSYmCg+P8gYRjN7tqrER6ZzSt53JDp8glU1UMsxezg
f5eIkEXWDw6N7PYLnhI7Bmg0tG1KMJyPDfmQ7rG2w/BoUUbOiL6LwEYfxiGkaCfevI2L5fYDuhej
lHXZtl6sU0eqL4/xrbdd3lgke/brBRYEy1a4wGiQ6MBTz3ele+9vpaVcqHltn6ix1oOCqPlMeOAu
nytOpCk3jEYuSx5uhP8nHn72X0n/qS8iu3mq36ly2mYec+EHKW4bIOj0VAwdV2JJHkmrSjhrCdBp
/y94HIu3YX7CtydGD29rP7Cjd5tphDVZW2Hqvkv1CrBS1OOj6bjfkGvn8JkQ66flQkOG8HBgjjKU
UOMIMfKdYUuX94jf6Ml9a8FwgHVUucK+v/EV++ATk3lil1NtorJHPhWDHiTVkS2qv6vIeZYY1YQW
IaxrX4BbfXgtJ1DVSkm5iQ0KezUrnHAWtxV4pQr+PxkW+1+yvHbYDNRa01Xy78dtaHLe+QAXyCnM
/+vQShhMkrz0ihAXw2+vO7+0FenfrxovWJvWfMmY/6usITIUSND3TH6aW3LK0nTTsjB6eCso/zn8
Ld9H5EUVAlt9jVvWDv53cyaFJmDVnsyD/6m62j7V5aspcwBjDDXS9zTrk9MWlCym2ryjEv7nYJZe
vDVRdu0ohwmTHDSaAncwTnATl1Ku8iXVxZLnehDLUeQBjkKzHqbDXumPCPo8m2R4pb52eENS5qX+
pDe+9tWevRnjUWJESY9hWwkO0CSiwk000qF4w3tUbjSNpuKdQ8t5jzRTHM0wDooUZanQL/NGpXpa
qSgF9dmfSbXBaa9KHhoM9zzOHRUGMEisJvCc93gmUoGpTi+QBzOwTwnP5tYLU0AVpWqbbsoPRtkA
4Av4178dd/Rr7irLRNmTBvpybENCGc90JPNT/CLlM18WU3BHeR1XhfrLpRi/2P0JoQhojX/LEHxB
vHf5gAqkXg7CVHe04WbTYWceJZ23gSImGufg3suWjwlnPvwO7H4oOB1AKYtZOiS7ipdtFuoXyi0y
pagG1kevIVeoHyprOUAvGwkL1SOOtF10kynjyGvd9+Dblb6lqDFuNhqKFcL++zAc6+S6BNZr/Cpu
HZI1gA6oiR65dP/4Dg2ATZBgQkfEhpHpKeMG3om0GxJ+M+VAkZjsTm+Oof37apyTDgNW8lZray7j
9X7iADyDYYnjaX+xbXtIiDCEgG3yGWth9KdK0eSsTY5licwDw6nyYTFwW3/cxch842UXGZdeBIPm
dLhdwt/NvfjSFR18TFry/lJ2gylzM2pxWs/ouO3L7gDkzWkixtBCUAxvISZl5zR89fdhL77j4G9V
B7m737uG8iE0Z6Y1Ak8+HDCNExNzSwkUdozk8VH31fBR+D539EmoRyoLJV73qt01FedRAA2cKWy7
6FVr0yXnj83pkDjnv7U9g0DJPlrCwqNfrSPvRKOfXdlX2y6t3LL7rjOhW11TVxXJaenbfnWqSRPw
d95EPHpp9pkEg2pjiAdGxxe5MqG1P6XJT6LASd9YS1TaPQinp46Ad36t//FwkJdil0Kzmcal4dGQ
cyxCdleNL7DuJmJNMW4be97jkbA/jKg+gFkOeNo3Ggd6k5vfbKH4HLLmwu21V1KNGtsZBch6nzii
IGo8JVlRIeMFWxccjAK6tzwGKwx7h0mgfQeklT/dmxAUE4EnQwoG3zENSoMqeq0z6/n/z1eOU7AB
+t/QYafCOKKbxEF5s1HfLiqeATYQfp5Bxy4ZOuUJgMV4+5OUATaky1MpDxHtSRcndfE/fYZ+UKOK
aPm1ihRog6/uHEAhF/XjkZwJkkY3nGj+SoRaI0MZsc12n47XyH5EhD4UOJwsT3M7UFbZS8ZKlpov
BlC/ZnYghRreedoX7hVe4v19NPg9R4X8tU+rJ+0d+Fxhw4iVyJH6YmEs34q0FFWfmS8TxZtAeTra
d65BOwL+Ex/5rDZelaHximFj8NbTuopSRFOkwx1W8UKuWRJKaJ8aIN6tzDMw23Wyfbg+6SbpG6Kc
4Fh34GNvVV0f/9gYxmTygJoZPb1KkpiRBxr4QodKgpYevKoovqXbv9QnyJMQQZ0FbZBBMAekx7du
sDDvjlpcKPuH4185+GaCAB/XgrT1tjsh1PLdH6AwJqUt8H574NumcaSPPSLJ6cmzf79JJ6MiLEif
8qm9i3retFzLc2xnLaUXcR2wU8SazMwf6agRdjfN9ebNF2e+gfDzwU2aw8Y0C9qUIjHWfI8wep3v
xbpNANruLCrFtVgDXj/LtQ9DLfQXwG4L/a/TLHhed7YP+BJxPMF5X9Mn5pTlZtevgTyGFWHlRVKO
Jhh3HKK3/V1kFwLXXisTWT8LXpT7ZXzKjBdQUr30WHXZcgdjdLDB1B+ex0IX/NPDkF/thQl6xmkK
1zBXTq72EV6MToajOxLJZX8VmkLy7HUSa5Y2JRU1V8lx2GDqUWFW6ZO0BQh9IzYqhg6RSTQmzZJK
I0laI5g26jxy05kZujrw7UO2QX4FEDPA6jGVoZswtHNPL+ShVKhjbwuHP2oM4ni5vXUz+XCOjMSN
ErGnAOIP3qFSOIhnKs+KrSsYdutYd7tTqmA/8wNHMgzUvtiwZt7SqoUMOubrbd4B6Qyu8Muki9IS
FtQORtCzQuE1+S0eoYCekM5RlBQmLblTSWXWU1kmljeCoEURqkN7J6MwdFqyCAkqaiM0QAz/cuAV
1/cnhbTASKFVFOAKi9HkyqTX8Ah+UfVm72bGwfC81RH/2nikQ74dZDsJCfPrbrmPVFmmiId4cUiN
uOCf+2uVACeV69F3VsFdrUKBsvlDNxYdZsv13k1+q99lmRupVx7IelqFevGx8tpd18kDpcw+pNWF
Xsomcf1efjIRqmjMKPO4uxb7P/gMxKu51GTeSMv4LR4JMrlhqdRuwebR3plCTI/aLRn0W4kWZfuX
Tyu9Vwbd5jCMY1ZuLu/rs1sA36g/VitOPioriaI1PPkG25W5ETPAXAR1xMBChNZiEP/rUAZIpQAb
jld5PWnaaMPn3n7tjG9HUKLhMdsjuvDU5BighY1UeYhxHxGpgP4OiODUEg0wlxTufJovy2PPrRkl
GC3rF3f6iWfMwwZO4QDa8cdT07JnoLNR21bABlnBtMve7rq+byjXoFktnB76YedkNp8gQ9KViYRi
HKw4ab0WABvjyGuOp42s0N0Nm03GPK1cDk8GuvIgGNXRU3BzGkGg9MLa3w9VmSfSNiQi6XCdtH+0
ZUIC/pl+Gj4rf3d6cfhnJapHwwoWFGKtFVYWq0WkRqYvALAB2K9J2Io9uZq9hl1aYVwPMpBtFJr3
JaOVJYx3uevZsKaeQtjbJkk5sje+KbX8cg7VOV3uh+Woz9yBxeN+DXQXZbsy/nWN5eun8XLrGWun
Ucv55KSe+/2bfiMVPtBmnPeZ1MyvPu5ea/CpMonItbv0AqRCiEQ6AnUYWGotlgIDq4VVIYDhtxQv
yLRMZyaZyrSkGbEatGAD8pkqNIEW9d3ECsi2F4wYkALG6VU72T1joAHY7TqYN2QdV2/us+yxMTY5
3ICrM1LxoHdOYvnUInJ8dU0o+aPGq+S2NwOEvW1n6YjsDKIQoUGq2436ozNz8dSjG595moN86vwU
GQBeWYu8ZpdbHz5lTyHyaHgi83HlLm+PCL0avMhqj1zo+TbeZ8W+7NIMiUsTXmuAQ2+UfFyY+Fj/
RCGoWKYC4sKBLfI63bzyOfL0Kiie07arFUWvHXsBDAov5WikfkAIOLNg4/Uee0IoK2hHoFKnW016
3EBN4/jeN2gWof98puAoISkxi25Zub0RDz3OppDrEU4tgFRFprwomMsAfrnYGZC7yt+qqSADCdlu
x4D7X4bwwEGHdgbqe/Zjmd5aAPwKYMzMhxvA5WTV6Tc6TN9hguT11Gg+Dqm46VHXA8A4BW4wtjDx
fhu608KvO9EaFc+sh4qdtdqHt6qe8X/VUCe6adtTQOrowp6bN9Dh91d7QRYoACcopajwf3ap8Xre
VQPBGvDMOEAfXGEcoipcysrSS+slYMPqJCRsorZb95pW/oW44rnlGe9Zjb8hTd20jEvRrQC4AFrn
0f6Xcshsdzyri5lArqYZR+xhCWFlHOCyrVhrcudbt7oRNdJ/HkrE0DxsYzhgHLTP+3w/guLlrKvx
+0AvneK2Cs0b217WbEX1kfbCJTk7WFLbn33GwabcSK69e4UBMms/KojnHpGj2ba6c7cbv1280DoM
JgTGnyF7nsXowYhSkbnp3ItMJpyfUKyuXtLBka8A1sVU+4D+DxBA3Ti4qaeo4y1o41IRWpwquxMD
fImF/OLfJWqjNkIV0n331t1gLTf504vmidpxY07l7t9qpg8HjnDwYo0l2SfKN9d/6aC63/LUjn1I
pSTG5AlgtQpA0nYDpO7/sWy5SdWB9gazy7Znz6J+KKttaj5xwWGhTTPjq0Kl2V5iyi1piNP7Zn5y
FiwulCaxjKLR+Vm2PXwJkILUv2TNQBtiO5E6eLy6vZU+tEc6nmmBDKsZSkZj6M8uNHTu12KIGAfc
LreENnmAIoQmoyXlpIQjkOGRl9aXL/zWi7+6vIlagDg+1RCKhd4FnJXClBj2nYpYq7uFgipMCmNt
SGHdSJlR6e818aqb9sci/2oTmX6L6zY7wOfAvItqVZDtIfIM77XFPsBoOmgy1ETKE3+EHPohIPRj
FtvAnDedF/XkcPcwZzOFj77iUCSlf7QyT/CccJtiPn1YohJDsAnBs/fjVoPGZ19EPxGGYUg8Ep+k
HDy22tLBFcOdt/FMa+AGmsm73xSgV34HeguD4DgU16DAnUUyCfu1gEXzDRrWKUlKc5ij39eB8Z2b
3ff3lwSifu8/Sw2nmxlo+PriO/ODlwTHVS27HiYEadbZbJ1QxbF4kGkZhLJX+RVUtP9vpLszEbd+
cpWlBxWZBk76YkyMVJkXUq8cwrH5Ztg0UwLRk27qrapveOBs2uziOh88iwt/04YhFgWH1RsnBZPn
RMWXyJwZQIjgchCzXQnWjoh4rcKKKm752Evqr4qCMZH55B8vmOYKty83uGtWb+6HzCQM/uXlRdLb
sM//XW/Ooe6QP1EqAIzgdn5WObO0s0M4DqDUMf/9JaWB3QVSxK5K+ecj+D+osm4UKOgwAulK6pKT
6AW0WTznN4XakkWvm0xKiJi+g8J9+pfznXhY3yoQ7xaY5iIlh27fCi7vlA1lMCBN8UwkISp43LzJ
LO//2rq/P6VBeTJxlaDiLPr05hi5ro9VE3zeXoH9P75oF/+8xLz3h/BgRaBhqwQ1b+7M7DRqw4VG
wfr6dU8hjkn+AeMDXPRfSLA28bzX7BevaHnfpI4XCcWVE+qm4Lm873o6HghDdtBiNuLY9B2gYirg
AZPhFWmrktSnRJH6ZDr2roea/HgS5XZjzUYPrHt69YWuwQXcbyIN7QobX6lvC8t9Jjf1sbIH6tk+
Gsbv49WlRNhIM+gJ1FxVAm2A6nP9dGGlnkMVwp4cHJcKEa/Px+UmK+8TvxygC2B38W2ysXX49vn4
4C9wm3AaHAdJp2Z6n+/2t+JKw7DGReyvNmyDt4EKQzcacNtdgVrFLEJZpxdWt+vpmdlv6RFWVgeI
NK9Sy1UMpGPFTCbGMppxAZwt81pYIeN50KlebHPZxmvu8rTi3LOBFXst7taL2vXinu4f3HozVYn5
9DKLmfXxV+kfxyTP+scD6N38yX+9llTphkQgEfcBjzzFilZZ8ffJM5oA2aT++lxptz6ow7PyF05E
j6hf+ehCHnfrrY2DoxfiucaZyZvd0wDsjCDIl6yQIdkM4ZzDzoblR/RG/SeEq1/83kxYjY2GVUK5
3d3DqlKCEiGHt0KzghG89eupA9FPJFcFIgdnc4eI122NRauxCkhYGODd+xU9N3bH2yq8KKG+ppn7
mYMn1NLFhmjAFZcngbemujg8xw3BcOe0koKDZN2kE6efAcxg+mmyrRgik5v3pUeYiMelbbQtw8IT
MX2Hxl0msyUG9lv4iH1naz1dIDG7k4mDF6/D/rfbXG5C9XTjPYu7oYwVyjzyvonSPJLnQ6bv8XUL
r2tfl/J9a8NOLwCZiYjScA5ygt0BZhcfigFylXvWIMoThyCHA2hTyco7ltY3TROgeH39zctCDE9E
JywEYMBTHu+PcTuF3UrNSPNJSG3t4XbykM73un+SUrwd1DH8m2Qs02owMsWNJxygPSxWfiMoHakh
DnvCcEwANJpkAzdlHKlJ4AlB5O4ZoL5kGdoGObRu0P0qLp937oacxNQWp/FvCbXOYrV6tmjtrCJ9
2Xf5T4qFuJwyc2H9NXtpTMWeZfzg15/tt9YcEMsFGHUt5F6KuYkjGAGQqumB1tkE/dZT/rqCRPs6
N5fL+3reek37ScIPWPHbBxykHdbm4fBqEEC2KqBuwq+TBZDVhpePkleoYLIesdP8L8Z412Vac4/T
cqXO1mONdlHRUz0wfo5ggHbjZ9PdW+ukXn8BZIyxAdU9eEVTuHq095inGq2ZNqk40yLxkvS7WLDo
FUzRADKVa1Bn2eZQa8U5XNAnpEXGrt6ckWzTEchGXtkt790OmJS4FrwfOrCAJXnOu5IoPMS0bLwM
+Q9jpRYZySw0TFcYKJVqP067ZDVt++CpuWrWtURy1nLM4snNfapWJML4aceILCVIO8GocRcStIjT
kBIO5WObgbbv73U5W3ry1IW5Xq60PaqsnUbCuc7B1/XspNdKpQBHmjQn59pnJWi2TIZD/9vSkUFT
8Mcn7UESdGAMSbFGWx8NjUR0tHgBQd6a1EJ2fAJ9ztN/NRTSY0WtPX7fE5xf1N8eyxQ8+XDY3DXU
yG8b8h3zHRWuMcoMoZss03cNrg7QrRe3vnMx/meFISkJksBLmBjBscscLq9mcsYZbAEKeVFgSvmI
z26ByvaRd2bDI9Yu3AX/RWZfUbcIhz6J8tw5bs+cPIzE+4EdloB0m18d4fICtVnlHIsreAOuark/
Ef0prGZbrhIMDAMeF6zv5lPillkQYB6scvCRfr5QH0oo85+vEMfCdDYSii37AujV1UexrfmIQXBT
lsWdnu/XVIZ+l9xHfcaSprDKtwCH0A2eqwRj2Yn08exec64J3Q9Q4akLSHt3FkTbQFm5HIk5lCkq
Ty9D5dLNfgoR36Xxn4l1QJ/fGDfn0VdgDl69731jP6wsSieISosU/TK2l185HVfw8Nq51bZbebOs
qrcpOe2wppVYHVilT/e/N4fd2ewqW6FgUXYlkZvBSk9XP76g4D58tAgL/DBAsW0m+TgCTli4Qex5
lkLfCeRUHiqiXKpuQ5f7oGZa/NcDo5aPGq1mKtDwQ7kGqPXPU8+8yosR3hUdhFjAeC1rM+A+OpVs
45O2vbxYoW2PkbZOdjO9/lBgN4bFSL0CljZZ0/V1cEnJNjq1ZCmWJlkgQfg7goQfX29iN62MsDmj
sPOxugQwdCru+Na3qt4bnDvoGEoMUubyjp4Qj2UESh4Nw12eJTgPEVbw+PT0VnOVNMpjggLj7JM7
3TUf6oxMfJ/0tOhSHyvjmWnxNEECPhBGfSAgWLijnbFVwxGxCbL0lDoh5/a636GL2ytRD/lOgzt1
ugFRYYSEysUiTdXhCX78Wa/SSKKb/mMEqzAxOZsBqqhKqpT40pZGugz957LLI8xNx2ZbjVqS3dM/
kcru1Nvtj9CX38bd71IHAa5Q79jPCEN4Cg4wCl0KNawwyrG4vqti+dmzp1Qe35OPE6hPc3yEsd5K
ALdDDJMsT6iOdfHQFFjEIpj9rNzxTnO3NHz9eaW5XYPvKA8UEjPZlOsznyIWPr0CMs9uah6eUkV6
JGX5hOvXIvZNQYZrKzeAeRHPq8zbOMTGawD3dmkghTADPdzX7jnTVoq8gkir2Lu/KgU/8+b64NMZ
lzt0dcLMScUaN1KJDJN+11Vv68FTovFPwrsvsOnonR6h8H7tfvhh3CnoaTDNgePDd80QYw058hzc
QEXdenP8zbbHJzOroxeqahj/4E1O/mPHSGL0lEVam3ZagQ6DTMu99wwoeQpOKggJNpFY/JUqkbdt
89/Tf0s2js+CFQGtLJf6BKdeTtUstp5xWsfGXnh0cfGPoYg/iff70LwWHG2qnGTGsdnYJPo3TPbx
8jVDVLFpDcOpHlyw771h2OdzeIiNbf9wxMLqh5bQgHMJL6uG+ZkW/Q4OkgYvoSLwFHAXuOqrfWOr
GbvdxHoDOu0oraInpO7Urk4mwLr8OvDxN3G0EM4VIKuyKmnQ2JkVh5AwhIRCK9xa5ClAPh94CAaN
MugSJVJf+yAmv5WixYQL6m0KjU4z0huemNIem0EtX7ZCAmed+6SqVnQXmGy3q690Bi68StkTKwNK
p7HwsODO6DrUPATLZfutmRPqAqk5HaJFvzqJXNfda8EFmg8C3AS7R7DkIrpO8v+x2Ad5zxqKPZ0S
fTaKrg9o7lJpcNS/vyxhbiN99WSyoebBICTMe1SUou0qRjTe6qKERIQ7EwSGYT9XtEGffb/CqxKH
oEdP5ZIbpjVanEqkwPUWsbgdLBnaHAWS5O5ZtP5jdn7GbSxCDNLLT80wKk6nSFNUmZqibZsWVs1P
9Y/gD6/h3YY31cWSkellXshFMdrE5XcyQspZAgMnlqDDlzjQBe67TQ7l79I42lbIB12kZpFg3ZL5
Iqwa6Yi7FFn2kCL7p3MhO/uHxsNW8lQlsys/8jyJ6uUsYr0QURe3DWY4mctA3kZ0rKRhnNYLu3ay
tb7JnUXBbvqq52yAPfb6x0Pkaf/F7IWQD2O+mK+795cGFq5yp19HVtpZoKwG1MNPKlkgfYXIP2tQ
dmr53ZqIOUpMojlIpvRCsUiE1X5P9cW3DUp5NHpomXa4hXQQp/r5ZRz+xabnNrYDbJjfKDGm8jTY
FtE7yuUR9RFvitQ2z6+iqAxEG+3rSrrnjEiQSEJhFK4Yu1a84P1JkloJHXlSxGmEIiagL14kfovU
IK9HnRPJlOrkQ8ESRpe+eXVGXTYkp399NdCjiWqGQ6RpR6w/uY9iMgvkg7KVi0puJIxdgavF2txa
TPLN62qfQkDlx9YF6koQ7PSkt6XwNG0+VEPl63srB2Zw/uxW8E8G4PX+h+29V0zQLTvY4T+wLIB2
Tl/QPYMNz3n95LOOkQmh9QClY98nB3nxYx1pPwvd+R6W/F6qikVDQmqufHHsDQouZjB8HFlWOkbl
0IwufIb1/2XzFm6LWTgA0AZd1eSLa2aluKxiKlJ9PrCJRFOW39HtAtvGxDUzCK+D96uojwdE+zCK
AQOuJoQyXztIFtAUu4UOZFl6GPa+fMlDgBHcvvGAPl6fbAJWp7c8ea2ITxic3mb0nVni7YJcaVyy
UGdNNUWBCraZJI4cHdt/wCeQ47AwN4aVJYjjvkc4P8hqVsZthrx1gb5On/k61TbaGSAhytJeexCk
FF4LXbumN1dKP3uUHR4BQYjb2LO7FuB9WCM5lTDZN/X3oxsBfjW7jBq8IFbHZdBGugbAwEg2G73m
LXs0mTPZxbAsDWN9EPEFtFm+l2ggHHtt2kvVaZ1bMa+t1waPAv1VQ+onBCYAKDH33o9Kyp2LlmL/
ybyCmIyApUKeyIQVj0dFqwfGaPGH76H6pxmPFedmTK0O1KGqzou2QIdsxt2GtuRw4Mmvg3VH9X5j
YzDjz+T+YhIi9qyNqSoiGfBUFJWXAE/NwPcGXsJwBZHGugYoiENyiKdtv2uaMK2LGVHEbetl3nkt
1lSm9sle0qy9x9hq1X9T2Gjf0yBRaNsjTR1tEI5MOJnwMScHA6hqg1XjueFVV5pEpWq1kYTIhQnw
dbaEV+ufLGfs4WrNFNv0k4HQmP5/BZIX2h461vcUJ7J+sbhDfy0aBnwthBHJJvdFlinrQzBBv3xM
7ta8t6Gnzz7E4BnKojlo7dIind2V5rFLVaQ2Tl85TiZ+Iz4a468BuUE5nB4x0y88gdR3JpKueNL7
Cg5OdYk5yD++bIXFcn80ChcMYDPm+Z1G3QftADwT4woyzP3fjNGDcTyOJWVrDL4OiDrD4juGWXSZ
4aMWt8kcQ/QGQR80S5xIpX1K0OHjeVrSDA3Gz789htRf/dmwmBxDU4BqREeta4vcf3cvP3Nm+oiU
b0+BfBx49aDSWDakuGghVroaycFiwJUX9RvGiBDOcHhvzGmulDKMQ8/blD7ZSGlaPrnpHPmR34S+
CnvbzkT94dUiu4SFzKmP92rVWU20u1W0M9PdjUY4UPTPWHqMITj+z5HRWavDJpAqmzI3EtBDGW+n
Ww9z0h7K2d2rnawKaHFedHdRdG9KQI0dSELh/yTLEp8prHegkENM9vE3r9dVAPD546fsXUWdp3a/
IdcqbgX+m3gh3Zh/E/wsC+Ejomz8u4IMFZ5H6xRZFtB3fA4PzB36Zt4WA5ldcRgau4NAYcJHbZlA
ePvzireD5HFIgwSArr3/k5oRpe40dk0Qzz2LA8dbk3NavyBZU3uK3XhAhGUsA3lVqcNLOADaJL4R
y3MJjXtCMvW+k0Cq5mOS2OuRm9qCKWVwpkc/li+XzQjl2ytWQ3hwP5JfpLyPQmweYskMpcrPl54P
7ou7UTmIOjDfrzNSn0kV3mhQgU2BJZ5bQ/swCIUaYnPO7QdZGsSCkMF27kIpNxtdu0307d/hoKCg
iFq4bb1f+m1X/2dJAZMZIAuQIcihi4rcMO9vW9kUKhDym6LldVEPyRIdqWOxGXIad/XFWrxDjw1W
G0N4yATVuxlDC/1hx/G1KXxZhfwgEAAbCs50jlAwRZ2N+5WcVMQZW+ut+eYpTmll5OvwVUK1POE7
QjbmQRRKzzu8iUsk3r9QGieewwEV75gLAN/BVUm7MLI4Q4PumI7tY/39gwk5WIFUXVSO2P+KKAsz
FtK422MkyOmTE/idDRy36kUB5vFP4/QwdfAQGelIvQzmz6H2s2xNHNKnK4ruS/Of5KuZTtiX0zO9
Yk2ZoDTIGg/x1c8M2kcLCNFdZChR6Op2/fhE3N7lmdg395pDL/p0Qtiwjo23Ndo3MXDbsMoBFLhZ
z3td9ph3rcxr+hZEwIoeQBDnrn4cfxcp5z/LeuJCA+zTxQ365i8zia7XNTNXNY7fLZSVcCJOSvSY
RopLixexV9ptwjYkBnJWKoDNcL38p6ktgvWMZDmskxz8EIpXkaycLonIdn0snSEK6tyZYn/zjl9Z
W433ltB3FCA6w1nLDEKo48uRw6wyBu5faHuc+7DsDjgsOp7RadPZTgHxTSn0AQVM307pFTCgWPL9
ZohpMeoLhW2tFgo9Raea3wr93vtvyqWTuilK/ixaUG6+NKJHioPZJ1mfaHfWTORQdO95d7pYozIn
Qmp12Rv1f8COsAWqiLtfQy+fbRnfST0Ynj4L8endqLGVSgoyvjFUguQgRLNjcq9q4jpaGbZ324hX
nZ3Rzo8sD5/7EWSt9s7JtwMAF/OJNRHJ6namIncD1t/goPyXYzZknXgsrZiqPPrgMYCe1tNUvQI2
UvuaQRmF5c2W5dF10AFFOKbmiR+uxaIp5IiX9qwuUBMJ1gyBs/KCmotoYBRrM4Kmf0yrhUoMi/3n
YLXW9tmoyqweSPkNBOTFhbXx7DsDY9Q7+7AdjQzlm22zJYd4LjATSrynqaQOqTcvIuVyZfPxXWPV
6rVhT+mx+79bAwwf0UieU1EAAqpe/pk7dKeSeihD7Aj57rVrAt2AZm5OOIP6u2IdidlySMGkMq0g
eKUuIjgbZ3nuyaAi6FFWflBoW7BPejTvOCtJEwwRbFYuUuGF6CWGHVEBKOx0O4XPgRo4ACdywD+x
Imk0RVgOOZHh0YeA6R5N7CPlnR7DrzeAu8ooCGD3+/jlZqXKEIc1yyulA99uxf/CGe99O+n/k61K
DB+S5zzu6LgoeULKhtPj6szpA4CVbTMQ7dzj6yD2RJkDztpXRVJnACnzmpU3oZogRltYK6nVRJEC
P+/uy5useD14zsLux0yAZIIb+YER7IwDGFCmDdNADZv29K4FULdcNl2bUqtowD5pgzCG4uv6HXCd
QT5PaHsYavpATkT3/WKLYrN8tZCcUPSppMqDrWUBGifi4EgapAH6gKMuqIhFg6PneM/TLolMpQEZ
fntpuDijKO6DSMze1W8JusDBQtPiuxthblNWn1SXQUUpLODoviCnorFCWx5j+6br7HrSfBHBRA5X
Mg4DcAN2dysArfPWdRch+yQKb8WzfVFZ1idFJE914dzmCeq38jt727E9yLfiqRJvIqv8XKkUqhB3
QSlWt90zkjqAPRjYaYYsRaDZxpbqyTfCuLJcf6i1qyjCqHS1ORkouEdxK6/uwzlFSpG4EnjvLS34
3uqxEcbjyZPurkuZ6H6orRqGQCHSbqKERO0GwKcecZBQHpSqdijZshN6fP7n+Jq+UbDLzaMwl4LC
drbsL8m05RDIHsF9jvCukjUAqKKN2RrE61kkFjwDC3Gg14ET6//WWw7RLUIdanqtIOMho8Ojf0eR
JUEPDwV40INbs5uznBANWli924x9++yeZWyNdkhuvGLS7N0xdILsPxZbn5URSvJK+TASssTy5h25
c0bSqMUFtJjevYom3o7nzIuq0OWZfQnIUT16yTG0ttBl7g/rVvXj4wd/rj/Jitj2P4IZTfWAo/ck
PBQ7c5UH6pmqlg1bdTKSRGOWEjnrjGK4HOJYQyRAnYlIUyJmttmWSWoy8rSi2NS5qjxByixC1cMh
Nuqyuz8keN7poTwUmqpVIFWhBrgEmuDEDUPBSnw9loWHdyTw3m88i8PTrtt2uxI49WKbxFBSGzUo
Yekg9qtrPuEN8bB6gId72XpbAJF9Di1j3lUHRdq3oYflIaf3GCemxyAvg6FKuHHL3wj53+TCXpzx
kp+uMkC6gTUdIEfauWPIQTq8iQwwsZaAxLE8JH+Of6Q2RZLW37Dsh3Ufyla4YAlUx5ZeJ6bsJNaJ
kd8tDSnG8P0y5KlXF8ZnP+XY5QvJR/QKXCGI2+qNtUGQ/GXBIFj9qzxF7dy/JTfu3pSeq9NIT1jq
Q8j9Jn+0g3X07cM4ktCb0GwBnDKpnIZgcQc+/rHP2R4xVbqoAQStxQLzkhCtfIOIIeefYbl5mRKh
sAyHSYl5svqnraMvTi9YPgqbUubEFx8xJij0o5jjjvYH9Jnu6tP2grWF3p0irlrtWrJsYaIkkWpr
7vdpNACnN4uTPv3XCZWRYud85p4XSuNFbBiqTYvIsfUeUwhfypJODIWbMRSs/LcMOr0b2jxSpPES
iWlKiiKaqT5mPg88dmtufvyrZywAKuyyN5Yas6Oc/MYy0+qxzY+b7fbCIzteMQkHdX/qEP9giwML
WdpzXTwP8zjP09VpjVU+sfX6IwpdRKFgfTXeYyi77WAQ1BpPyrhp2a1pfAmU1rprQw/3su8pIl+o
CuE9FN8uMVA+qI59rtID6uoCDS6GH869ojfG2T5OUf91Mgy6HJmKtNa2t6KKTw0STr14nFyVggTJ
SYccX2tCGyGo0P+6PR/ZkyYRdfuzlU8fkiuWw7OaTLWr43O3EBtu/jxhikIHrvuSXpTz0JlJpFgF
y3kbYefzm1FruNlFa970/c0Ijqd/UHDQzWOnK4T+/CLCRZ1PEzrufk56KAkTPWCSMkf35pu/ztGU
bLAuAcijmi8z50kV+rjswqrGES0dKxO62a3yUHS4LPjD9SjBtbLOpxqPlp2GRVcY3CEtKT5L8VWP
jiNlORcG8UwH7Ba6BNF5wlVA22xuKNdJalWrFuRL34r0Rh+r79vUtIe3nrW3zWwgHoxOHwtzTGaH
etUTEQzRoN3/fYg57/L2bZAEt/fNvGr7zszowj3RzC+eKDROBjF1chInGTNVYbMYLBvy6mttEQE4
wKyFNjF8dIZX7LNSi1AFQDl6l4yeLV4VIr7Mr06/qPwuYwm/X8ofd7ZlxEIUNYPc2tcZyEPcPEwG
29b6zwtPkTPKjUjzNimCV4vxZdxbSiaHGqhxAE1vdFW0yPYB+Tc9sZ6bTdcxXNTUuBGOGgMZek8i
UG/a9/ZKBrWB4DOdpfU/ihsczRkXgcK2odhiSWo0xNkSDvR2UnlDyn6W+VBQPZtGUuf7f1rgDVPa
bLcr+H1gUriPHR0ybTcTw2Jjuwo5Zp0gBWsV4dknNmASnEt8eV2mJJ6U9ZznppJcsRNDZA5pHM+C
MjMLbegFFx/vJnRwXL1cj4taWAfTt450fsMZrN2fldUzaobeT0hjAgu8Xvh6YygtBxUUfIbHV6ey
rJ9/VJ7MMEPt5No1DwpOAz0dl1v0FBHaD1magkk6qxqFGkM/oLkInpUwuFzsqe+7WWdWzVqDDZ3i
MwzTTGV5Rd/3wI80ioyw8xXmjkoSjPeTIOT/RipQbreUp8PD6lqnKt2qhGxYSre8bXNmDHz3rlfO
yLpvcNCwr5jVY9Yf2zxVHFIs4xq/M6AacGUrQX3vrPqEKRdYLmEErfVKpwS3/IpbtaivsyaSl3Sc
WO1U8DzNrM2e6ZC88Fv3tl940Wge0bjSBHunaEr3FggAvjAHFG3eMVWWUPxrlCu64uKwN9SVQWu7
ghV5Ck2ZMgl2pobldeqj2PRpKlFTAAA6GiGVrQt4lyAx2e/CDjJ5btkTDfqOTznDKdOOKgAJDyyg
n3BpGuQxH4ZcNYXgMwYxrO4SP1lhh0lEJnN2ypndMbxMgmPrWKQh1fne8nMN7qRysCqjUoYbqQQf
JZk+mAj25EY9NNJXYD7DjSC4kXW6XR0MDQdl4g866p0vndqqOwuTW6p9Fga/x1r1mocrMvgyD4Zz
WQD6q7k+2vNNO16MM+z9HY8KvYlivdarypzODiXuy9TvKepZqxltxcSxmOEvIa9iPKYkTppZfNvk
sO9buCEF81AKi/kDt2rDk+cZQufggWDRsR2QC5SHsiwxghCBmqNPQpQIh1w1+lfNw3THwmhhZ2yr
RGsnB1VMO1JbYQHk7lfdoClSWSs/PvKebYbZIIABFRyKJzP1ZA2voANGD0OGatAjc9zuGimTZTgg
sQ6XYfUNSweGdt00R3IkM6mGwrtJcvqOkErYOu+zmqVGN0R9Z/gDcsCDJAX5Ia5/g+4MpS0aNKmH
86ULJ0wX0nqTv1Rkh9eoyX2JQiD/hLGVnLuwXqsv+5HG7Oqz4ewie6xwv49U6clbCwlagtFJa7Ad
z3VmNYyM0EOS86rGSL4WW6MwW6UpshRZEvjRox49pXsSpKjkvUFHS0sJcBa3A6YgFQ2qjkJODCqt
o4DythKe0/1kuTTrWNggWhlIpJ/YpCTJ7TO2OnldJfQAYgz3BNIqtIu0/NszJNGUYi4Sd+I+3V2r
fnaF2t2o+ZYH9nWrWVHV1Qpk1/05HqFuaG7J/ZbCaapSHEnyGY2GblN5csUOuAE/0zIHDcYsXIkM
d4yA08pFRcUzix28Od7E1N0f9EV9ULcfAdNKZDjtCLU2ehyQuORBq5XyIzairhsgJsN+QFzODLnp
mUhQ5sXA/58zCQh4nhhKBhD1S6HFa1KqQlNDj4sWMu+UTOcXnf4sfKfEYudRsfUbJNnlONfOhoQr
wZcskCjtP0pVPFt8tAT1NYICAKhypBoOVVwdzyzQWW7End3AOrP11Cy1znCYl+liEYU0w/w8kJk+
wK6b8uH0KAs5qxjO25GqJwHcgPkbe3IaMHf7wxz5RBIewXchqX1ZGa+zcJBm/RQ1MNSEimq6rI0Q
wIUbplsueA88kJqm1yInvAkSoa+sRBCaKJHM1EMFxittAj8AuKBT8ZjnynaWYi8mtg/bMqzGUHlQ
kVNvN3/KU994crtlWcu0ZD5u/+Yf5afQoUuGzZpedygSLHg45Qu2RbUNokij3M3du2Y0csSNPf65
MoNryeXyIpTj/U+LzElQIg8P+Zcgzz+jB2taCtEFHjdBXzPGl0p11ArOxgnfa9a4DrghcNLoctHj
NVNgf56Qq/+0RfkVTO8ZAz9eiveQU2J715qppz2IVv5zXwnK6YUpN+EyUq0ftFcK9c4f2aHa8eKo
VxQc81Q4JqdFhtEl8dtK2QPi5e7apO/gBGtAC6n2h6r4UrB0un5rTxmsn81Al7HJHbK7SrjQvu89
4m4ug86fuKZGR/AD318E7I8WAhjOv0bWhPK5E6MIKtdGKbXA+ROG96bAFnDJQT1SLNj0I5yZ30/O
7DBznnNr6Ts8VEzlZkLXL5HEJEMIxRacsARqVDYJR3cNQ66JU5sZfhhv6S0ZuY1eZy8fTljliFE8
XumRTF/XT2p2CW/bPbZK6yjMHTHuKMroaDNrT5F3DSPHUlwsCBHuVtfMpOo9r+y8rRWSw75t/FTV
0h91JEGKynXgwpIni/oz0BwtKxvhUCoax30X846/vBHDd5R+Zn+UBjxUL2HQb253hnHxugpwMuuP
z0CgljjRICCPxDdlNSLV30Rl+HCGE2nZMSQQVogI2d+Hb4xBVTVWfLxalqytVgx9kjrmwXQEt4Z2
Ldq+hkZ+EKv/yvSLLtsnwdgwJ3KdZiIK/6NPyM9DcDBo7/g7OMwpLsVYGZKDRxbe0Xemma8Vy3fn
hFrYhcj1E9x2PNRa2tM1IGXV8YKRmpJeGIFgbTEmOo3epuQ8/ak5yyuDTB6Xqt4rBs4SC/HRHkob
hyNxjSwYFmh+f24uh5hVlJR5whn7T4x1BNPiF6gWd14t1q6n9o5u90ZHNPUxbpe2N7k6XdvS56mN
JvSZq+7PhG5+jNlDVVnnXuMnRvzHatl18E87eOzg/qmstJ3/SIAawqeosmHausNEo8ANQUJMKJeh
xlNhKqLrhkJXiZ24gy3zBZY+79IALsJDnFs17n2LWRBRkSluFlFmP0DJIOc4KAY9qGwKFXx10RLH
UvnJUzYMh2Pe/ZCLvgsw6XpQ+CjCc2/3c7hHUUqgRH//KA7dUbGZ1JMM+pighG0ZVWZesH7RBFP3
cvgd77R4V6cbq+jfIY4JfxhlqrZrd0TKFRcPrA5Kgrm7oK0mjPER1ePeY4qXRg3QvJTs4sOf0gPz
9SgZSQWeR5wtl4w09AhvNH9iGZAO1JKrmp6qsJsMjuKAme5AQ3SjAwau/GR/zgMxHZCZh4K7DNMT
HazY0GxnIuqQAJEHArZ09bNv9G3OOzlDWNnCl5hiMe+gpok8LwRYzddXUA/xa5ozJ50DKZrnTxiZ
oSFLbILPSr4vWuFJSqv4ULSHSIMhbAfEo1EOocprYq3laK/Kot/Z6KB8SPLS5UVwpQmMZPYhP2ek
YFDcoqEGP50ETFEGH+DZAqanh9DVvCntUMwTHhKJfB6BhVSQ1pD7XTAX+eWVWz15kAShePFK66ik
sp6Rhlj5fSbw/hki+Au1ZSMo4y4T/i+kMAw8JDCs37GDZ8oimht07AVfiI+bc4R/AaJ9BCxHwV+v
2gX4JaVhVT3FXl9OyBEIsq3H4Lzko5JqtnFO4Jc5MDmnU7M7VYBR4K+d80mUaWeGPzfJ0neBClrn
Cm8yyzQH/eUw+erj83EdScamjDF3Mrw69FCwPUH1Urv25V6a5fWn/OTrJkscM4Eu7Lx6+N7BvZ6I
VCirNdpsZPQuc7Nuug87fGwE5aU0GdcmvYb5vl8nkqtoPDaD6D9Tup9obrJQKtXDhm66FldO7l/H
Y+XeISw31rofNajNCQd1G3EUK0L4j1I4nnRnlU767t/wx+kQZwPbY7YpJfSroz9IE9zFYFdXSxGM
q18NRFL3zfTj6Td1TBLjbWK26pIwYwD1MNvkP4iHbAo3Vhdq+rv0a/AAbQhcgV7Y1LPhh/+1oFDQ
kXzoDJrzwt01TbXWcvD/VFDhZVMwqO0wDCWIglZGU9ikiu15a3JaabYu1URx2lEONJX4EsspNfVG
NDhw2OXH2+Q/n6NeC6vmPn3T9UiYZBYdFqJmUM+nCKGy6QyMvsKtlwt777bgl0ORp2blp3YsILvG
ZPbjeBRw2ef2nG1553w7cFBF7cf+nOx/AmzPpPDeqttKtWgCEGBX42xcaK2ReoTh/SZraQ0wNdkd
XAYVwQM4cAqsoy5m3o3gsyY1tfsEdFThEnElx8ezdLqFMPCYaW8w+055rFtSKVWta+bMhFSthoQF
QgvXKx1jtlZaxNiEwXq0xXOAw8Z6YjXlw7ieIAO1kIsVaQWEfSoXw3lQ/ZFVkSROOygQ+mF9HpoI
68syZ3r5tQb50N82NyxEAiGCVyhGMgJDvSeBEnLanQnvLYeUmydAreInIpLirWikcT8nHV8wkTDr
hWIxoVMOFdPDITcqiXsy8eY4meULw4fn/2kByBCcLjUatSbi5yKxLkrXTUGXyl/5mWrPFUmjs+vy
4z9hYMrAaKSm4ZkJYH00IagOn1jAKd2Y5h+Bc8Kz6vvzxAOWBqioOgGx6AG778eJqx6IDilRXIUt
7rQ8LZ3iG2gDQ1dCN4NWDy+U3jHRVtDnVQwQ8qz3EUqZPXJ/TT7viK93DziywTrt5xBkCwVVEo9A
Bz58BLOx4eZi3z+3NzO+tanre9VC5WPE97ZAv60nTv95Ayn1pxSY3oQsBZ3HjMe7nkRK1DPrzKFk
EKIupuU7DN7HBKcbiniiXbNVx7hF++kNbQXjuU8V+x2CJp6Tcp8DGZ+CXE6Siniamgo5HjFWy5cC
2KIuqKFIZ2r+qFOtgPYw5OwYRp0K5DILAt7sdouDKVPjO2mGno18m0KYML9AndgazF+sn+onaBPT
snN6sO5KHlvmGe19F+/0t55WOJmXABhIwcnqESz5LvTzArNJjW6TZtXBC+XedZ1p0eVHCtCgE+cj
nNrwn6GTpNbZ+99z+9newHJHxmm/PTzYFW8k+mR1UbfS3M/afUexLjbbfPD7ceyG+XdjZxuzhEyH
BBhFBrfmK/sF3bk66D2H+T6WqMqWP+9u1FWCbqTSpzaDzGjnQBZ7vWC0WeXDZ/OfxXjNvWAKn7P6
03IOCm6m2cr0ERUCd6wWFF9byMTZUSctIfX/afvLKHUPquXonYHkNL2bHk3oFyRpC4ElMkeLttNu
3YmQgmESAVSHYQig9tmsR/e3bJeSmWhVpSrgcP/KVblalOwkUBGWDRcyELX0oJ6CS5UhkUeS6GbQ
6VX5m8RnbJRE+QLHqm0DZ3jub1WVJHEyxmiVfSbuveASrqAnC7/b1OKX2Hd3lCmeYyBAMDdCNhwq
yfgriLi6QXo7fW2xtGdKb++o5stH/b6ShTSvtzCFSAwoKc9HtU1zKfeC1s14A5N2D35gyDfojyfs
3B6fuWKcmSFti3c/o45WQBKzOxw6q6wScEfQqdO9mm27jMfQf0A1hxuUhIrQs4WGubsfJTYglwHd
tzT9z3NxK+jqNirk9geQ/WUQ+ZJJ8P1Y9WK+ZPFX9Kg3Uz5Z7IFk7LgVRWTbmMtKolo2pmh8ixjk
G5hjsN5ysohkKAoM9F+w6gFS3byNXqzSyISDhaYzw19wxpT5GToq57A8wF6nWvPBUDHhj7v0u4DC
TZYY/2qr2T9BJX6tT2wfN0NyDCxF5EfnMXYOTJ8jMDjL07lgSi7FBQ7XY1q31v0ONuxWbGTb3eUJ
3MTRKMRpdBVIWNyO52cZ1R0N7ZWOJ8nCBFhkwToyBTdjsHCEBC+uTTX722HYXcBfY3znv7yWnENf
Wbh7laamh+ryRHu/jquPa3FmZFz0SxEvJmnIwgs7CWRKvjKQYhaLkvVX+oJXZwzrDKwVuoJ3gtbZ
1YY8ODqTurwhYVchBRfiGnupwEK3Na+hdGcbdfZyd7Jxp2HYDhh/8heO9MiJrmsG7HmEZPpA9lGe
u/NGTZU72YPqMiPRszx881jP3igeVXExED/rtnE07S3ae6Ngp1XACYvymwpv/fuRJA9VHh+g6wMH
Irbqg/6W07a+/bFRavFVEWHmm4SwEkGOLIxTl08hY6v/EqXut2Jr4rljO1rchQjfMyBO9wpTebLn
S8b0jz3CIt9NJn0/lhfS4oxgR6iEFA9KBGEj2SDjvkbT3bJtaIKMOdyKy0Wx4Hk6tI+iPAUzg5Fq
rStDPl2lP5WLOD6lG0Vy1DFmTTgAYXObRWQOMYqOpKp4z6Sy4RyVv43ktziUyG4Eh8LECZ3I13VQ
T0VE61sRb29UgXyopNJuYSUI7RHH5XQw1zW56ubpHXJrxXXdvDJeW5wTihXOx6muQdsmak3XCcoo
3Ie7/XOVk5EdAAQ7nsttV/9HyZIJphjWHD9ZRBlVIbVvhDPv2Xfb7vq5Az2i84ajXQuUW2D+fvMG
7Yxy10B4t/FIhmPGD6EM7rujvUzk1A1KJ9FJ3TMbbRt8RdB5gwP1as/Cvg8jn0vU5TKV5XCbPeNE
vdmzx/yla11G+ps5hLvHserVeWn/jeb+njhEVuyC9MbrDTXSPSWQp1un0XQ+cjZDu/MeQTj5OQ3O
Xb+hgniZiWU1RWfHmnnkDb9mbsp2+rErnp4O5+Vvq1IcF70yTjvEyDijVp5aEF5Ox7DHrXmruKgK
al6EI3MrIp2/dMldgxzvlDwIc/i50qRZ+ZYtBHPG8cJ2jh+4+r2G7ApMkY9R1q1I9LHyf4RWxCzx
eixIkMrupmPqZWjxWAZEFZYopYt9+HQurZnyhcxvf+3GC/K55dWjTTRFTevWPF6PlLJ3GhgpVbq3
6rNIBG1hxxWxxODG2CDRrs2iWg9Qgeshcq8x0zhaqyvwxtwpnMzRVWizqbCTDi3C5/cPbDxYVeEI
dpSMzuYD1ZraS0Ju7/LmXlqKNpsTaoB76mJ6438NAgZFpBTO9hW0nlsrrIv9E6uDku54h+uqiqpK
OgMTb/OCW1xss4P7kKOZq4Xr8WcR8RzGIzK+41SR8ZEliHQetVEKHc2OkbLtWnwBVgj6ed3niUNJ
+r+tT3kMimR2vXnAbiDwHRfbKsesxDqoyHbTyZ+E04mfZ1Lgr+/ssQEIDBlGUI1tggmZQzvtkOwg
gxhsogDd1lwswLNbMT8s3p5dP5/HpzZpH1ww+g/r1Bw60i1TDJ5wntkyfO0uSOKzDDLHhmqV1w0t
/LY023D0yRIAfs/T6Zb9BBKmjnylmZMO1cHx4+CcXXFaxgGKxibotqZ/M4eAm2E9FHuHYE+MaM1O
PkuvvDF8+3SNQimHJZnx/vWExS2hUHneW/GoAzqIizs2K15oHPPzVRYg37/HnX5BOOBgP6nayAot
GKx1tPGe8UNsnVoaD7mEzIvAdwWAje5cx3slHI2Y8VDENJ9NqzxNkUZcVZ5kBdPzCkL+zW+S6sQJ
STjHMTM6fxaXvEWwlKcmX2QF+0vkrIYh0ztd+fMCk9cj3j47Zyj/NNJmrBwGrQIDkjIPyS8qtLEs
opeM1PZa5Esyqy0E9ehj6fmTGjM5dFHtFcssTllbSLco6XR0hPfS8V/+THf0+KZdRKrogJeWQ+0z
Y30VL2bp9Gb50sOdTOckhk+fgxNwNKcY4DnFMG5nX6f70phFHOxK0W6M2MeDDPlMtV+lVfHWRJHf
TeYj5CXw/MVCnlti/F631dQoEb52e9PN2LS6GpFRj10bXwBkLv0qIhhQT6OHu/bwz64RPKU8UAPR
+fGqGK0bDfaqblnE4OP0I+26lsxpBYHM/NS08Lvg2ZPzym4DLJEZguuDNxIzeyWFYN2lVF4/Bd9c
qlD9J+GiFXPj947CIANUMb6ImwMTYE7jPjxH0xjEeTxNdL7FS+DopTr2jZOi8erzO/4m/umLFLhY
djor79RMX9qm3nNH303Q8pJHu1tMPC+tBqcaJeV03/jpkp6HATgThm8XDIxiLQhcUI+/4v0GBbKu
ZIx7HX3cLJ1o7mcnXS3RG3nKpNo0gz3JUg6vPA8Fg7lOnFFBZVPTFDxyHaWHDc6s5ru9izbl9Hzv
GyFtKMsfi1D4Qc1Cfu0/DObPESjGDc5FT9r4nXpxsJPoZy2yu6tzogTgGYZQ4IAsv09GTUdE/j9M
ljrGbPVhCjK0651WWI6JlJUw56FRJORDNHaFt67bCxzy+DcXHHWvvFoEv+LEuVDSMSjE9+VLktVo
zw8GdIq3AA4xlQKWVm4hCNdOMlMPxXh5PqJBTOTWLiNWgs9im/tVMQ3XYLKxPRel5qhNctt7lXNL
C1TjOc3CDIDcPaOxr1f3rxAIj20Y/hqHa3Bxs3Reng8KgLTSzAhtKFTNiVGvCg9im40mQsGJH8jU
v48Q0TnmfOv5EkrjWcac+A+jRkkfexbhxf8hAreGJfdiL5GLespQPLywIIPEpe4jjYfQvsEm5RhY
gGXIUCT4bNYQRwpV3c8Tl5boeCnotVZHusv55YOiuBbtbuiGaGw+YFe+/cELmrMZ3Mu7cYkgVZz4
Qpja2RLvt8G3AjZlEPo2WaQL+y7HmOEGtsPv2omCC/yRPousRTj4SAw2HLHV+c9p92kT1q65ANBC
LQniOdVvuxLroDPEzW2ci8gnmfDHJZyl7pHRCwQcnHqV3EeOxHXyrxWCp/O8nsFr/TIo+odhZpeN
4TdtdlQg+N5rL3KIRvIqjS3oSoRJgBj14uAi7dbO9O9DP+f9w8ZSD8/A/q2fWYiKh9NfFDzXQgck
wdIaoIlwYtseefBihyRLdgchTmo1eO8EYI5KQsmq+f1OGaLFa5lEJnFJEtGYQhRMjV6ZSoiHLbQe
UGA7O2wdSP6oZMtNwOe9mSuwxqWLQDgJd7puUNUmLkNhBLM6kk/sgpQeDFVwgNwFkzk/9uMDZkOV
aUHRSyNh+FKvhbkm4S7FR0xnibL8gtuE1jXCARit6HVZdhmK4c8jaJda6wuYTw6L1ESaYEE5kgie
YXhcGcW+xP97dlkL9reV8UnMMosV6AuvcPuWwG+HoGl/UsvbNdlAEf5SyNGlHXFmDAUoYiSanGBd
kpbdRgNo8BsrueltBpV0Xp4XotbN1SukSZ9YvP0VZmq7lixoV/uYrtt+Zse+ocB0AsvRuw3wuVXe
xb3pX5DrU3Dq10Vs62j5d90xNK94OH+4sOxPPtIhA74kkJyt7hp8c4m2vF6rHkEQB8AT68Jq8074
+ulMAmQNXNh9mTMhBiHUNizGxhmM2eHc0tw9pxHy2XQo/y7+ZODIQerm6XSvEqLnCJuDG4pwRJ/J
du4EoRwn3XAS5rL/oRe9kUFWWc/ZV/sKmTrtZYSLyJ5nU2JO5tGawpX9SlHFzomKxrUWb9gjJH+7
C3nkZiyOe5SZztyRv8+Ip/oJJi0OHiHV8GWiDix2L/wQVRx2OzFRVU0VWVmKPJBDhH79qH3ov03L
JhkJz8rPNzZQW9XPBCwoDGUaeNKLBXxp21+OM5VSyx2k6DcVfCXwSjmI0BW1r496/XD63BigV9wh
XGoRXNajbOY2n2SSu3JQJ+4njWqNG12/bDpwMcfAT4p+7IAI55IHT6VUufINlQSa2CqUV1fTpbMs
VRaWTI7+q/dQq+PU+cNsB4qTeIz6hAWdRgXTvHBJ/GUodrnLfjOQBZEKWed6dTWNKtqQ99L44a47
oMgjTFPA1njJzNHb/rKiC7l0i6CqQaSKx87/0Fpbey8xk20iZId75DppntxooJFLB0eFQtJUct7w
+4nQXiF03ab/sMvTiB/yRKkXK2/O2sgOzF8d8JEOydygaPt6+qOGYMM7hRXI+7HIY0EgqWp/mjDN
EaVSV2GwejM/ACUXalXkkTVFdSbtF1S/P0roznYr6QaDECoCd3P+Umwa2CrIM08RnOeVIKERZmL1
FFn05CfjMVqKNdO8EXL3vIhAT0b86bt1Pz2Bk6W0bO3nPQIvfCHhQ4vjQyiij1j2K/zysozUMpLU
+ZynP32jqR1OHcCVatvJCQ8Kfqf1jqx7XKmaJgk2oIa/mAevoHOCXYmmOzPGBm637R2Q1RSWjKQm
ICC0C3LBFrPjYDlnxMb7/t7ODBvZkbB1lK81ldxL/RPP/10+n2tNgqRilLBo5XmAV+sNdQ5Uue2C
nd5hVyI/I0d3qkZWkrlLnTccXCRvv5j6Hksyr6S16I9wjo/seMSJI2EmlcWyLKpPZoA6X7ge4FH8
uVO73yjDSfH4ClCQp8kxikwdGc9TU0Kgj/jjik9AioSQqZ3iikYM6sLnPzuXm9MnAoYy6XTX3HSD
DMDCn+12V9zrD+T1Yx9zzx8MtddJbNpQhztqxq9pQiinYyBMmY/xi0DkAIfENnKvsxStl2Iu0vlJ
s6R9DQRr/PRaDoE2wwCdAw37B8NKM0jYFHhW04SJ7HICQRzDaGcpCf8Xy4FlAR8ZX02Oid98L2ge
h9pVEc6v+3nqWtfeN24mC0v6AkoMYuHoDvW/5A6yhECNdwPUFRkAF/vklV2gN3RjozrPMeMHfU8T
P8vFOKzC9HuTdqfzRk/Jx0h6ooX5R1mAInu/esSDzLelzPvE2oz+akWHj71jJLatbyo50YbXpHJJ
TPAATN5ApcOtV6Dsz46reWDmMKFaSDW2DUqIcrOrO92rNjo6HvqYOTqwOgbkPztUUdCLMbkxWiLJ
MxFydHd+i2T8815N1ma5HAXyjfx3Bq0400VRxYNrpy3UphjrsMkW6o3tIY3es5AaqB11xO7qVfGZ
ET1lJG3M1vT6rOECsYFiiW4BO0hFnvxB6wTDW/ka3Xwi9YbjOv2wYo1XqrT5u3TdzJMtaRQmWCSW
s0rTGpoMDRggmZVEZQ4YFA089QPM9b6Z/POQ4Jin8Je3iCdxnRNZxJxyo74IzhGD7PsD/TJlNavT
mdJI3JFsRa84nfKdhTd8si8FM1D4AztPBToVMYjxVOlRzQGm7/BtDZ76PYi5XfSoWtWO8nQVBrdq
hMGqeGflCdpQGOrjd4LVE4aCSUr3g/NFJUacdnHdJJz2O9OyX7yVqX43HfKCr42NeBX2Z8G5bLK6
fKdqReQyM5NkMxmBxXZLVQrLlg/LISUaIaauEUVyarQNDBfiZTTXz/+x8tXkDuxXaANJrgd5h19w
C4zhkSKJpZ9uhR2xlDpj5d6Cddn9xdatoyZ/l1GZbhPMhXkA70YCqycmRuY6krAVUV1FdWiWCENk
yN8c5eYfufM1Mu/nrxVuPIUNP5nTBbVz+B9p196khhcf2RTJKnbWjbYlQFJgHRN1obzckU9Tb46w
UXNWmDgdrxsCbUeShWVIvOZQpubfLsxLQv83DWxhGPdg9O9LxkTR1B89YfpUm4vQfHDPwszOWZnW
NF9j0DVOrY3HX+UXb7GOnuj1lR4cKrxAVl0NBTKFn15n1JnjUBfrJxIk0aYTBQ9jqAcUGuL7rDS4
WDKcytVrWWEzw/GlaguvyID36OalDPtiW5OFsiV7dsogkLespLaV0jmBxDw5xy8nG+ZUieNC5FSe
vfILo1rb7hTyWAPsIwg+ejRRLQ+S+IJxPHjl6HHBqYZ6cEGBN6RO97tDHP0RVH2ooQx2g/eixKdF
z7fpJ3mb1OeOte9YrxKcaMCnV9m9k5EmZLlH8yJI/g05GNgOpA3XPF9ReTxW2OrXH3TnUKZvXQ3t
M3TqVeqH4tmOd0w0cgktNFU/phLMOFb2Q9wmAsDA4Hf/Cd3sZsZVhnIo1t2xD8HS0whclaBPFvsL
HnBP5PL+cOiZRv/ZWuoe5Kl7xEjoiImDHcSoP9HjgGJ9k8se2puH02VOsF8eF2yp52d8iRwZP0Ld
joqpmLkagD0Q2npX22qP8qgn7aOwDRV9lAnIrxqFDfZHUlYSjc/q9FrIAqtBXFlMrh+2QTFHAVFE
obB8u3uznb5C/KtS4249Y735bsBtyKROgP1nnwERPWXuQIbgaOQxpN3KSbCi8Ty6GYKUDq2TtQPT
CEqmvrL1MsEGpskgO4+uXjWxtSSMC00cHPGJzcPGHt6p6/IMclkirjjIBrj+46+7jyea6cjfYoBQ
GrOZz4AwRO2sJsGLJnVzVx2Eums1vQCLz+zA2AJoJ+q7u/Ik2v2bX4aYers93NntmyLSQ8GOCGoT
9Q058BIMASK3PiH03Cs2giqZORSKoCabXtzIM4sHHEsH6Jvp5FrhaHu11AwULNP0LVYpclRWGSW7
UFR1Abgkp6NBw9HPjIOQm3ohroAaNSNMI7+Lsf7KOi8nXtMSUiKXwLI3ttHKJMU9XMAaUqv2IDki
Xfj1UlvdeslWb8yBUfMPP4o0rpftCgdMOG+x2Xg2DPNzUUXSLLcukLEyxFufHR6dSxeO+GPJLUfO
KouwAKgK3ekS8yn1PA8AWCI6HT6U2jK6yWrj+F1rX6MUxEgGPDMlKUFP4sa1wOrOoSGvEhqzZYV3
8/PureN3ASEj2Lb5tiflYaGNTWKmhz85E7qfunQ7E1/TIRxjBvZtne4rfQt8eLF4dRmZxeTEcOjj
RrUiO4LPNJV21ugf/1W2mix3Rx4w+FeRYG986n4lPCxwWNJ3ix/Nzm0McXhvrRCntvp1N12iX/Vb
D8+gEM2YF0Nrpb/bJQc6b7mGMbS8I3htQFSkTNUOUPXrhjJ+QrV05J/XmxRSyDoeIeIbmUOOY9vG
zZ7O8wh4LVrg8Kvn0+O5k1CIJ/tqeG2T7YjpDbN1s+lu47axh3G/KbK7qZREDOSgJsVKXA7Fj+Av
eC03OT5xYXDbHQR+3MziwvUnZOcTpNTyFzaCY2noo8QDNnTlEGtgQRFeOMknTf8vEaiv6tmploSt
rev56//+kqzEjCCmfe1JSELZMFV0RnocVfpbx0thw6GXRKpLiY4q8Dk4v+2uV1KK2+Y4gn7WBgMQ
takZowFKcITZfZPJtdVUai8Zo8zTsZANfD938cgkcK/ng4JI3BC9FhTteUy9SlvqeGzyjP9ZDTA1
V4nIHsQiGVmONJi2LcQEXC16fafxOHDqfvBsml1nnZU4pRRMcbFmSSiu1Ggk2O2ztfBpzEUagiPL
FcZh3LWUo2si5xN1cIzEWJqslaL7IHcE5N533v3T3JUAGzTX33CoTidc9T606pqrXF/YpsFwY3x1
fs8v5HJVi0TvtmI7CSsfebmrmb+remr87wOS2RUxj1o7OWUhmhiFltN9wm0He28G5DYkl3EpeOIo
cNuTiS3FwSnxBgMTtM+t3Qns1CY6yr8WIbOCWTllP6eUNp/a4x81SLobUWXpUtcAbYvHNQrbyh3V
zf7Xxv1w5QXQUkXtzmNotyszgjbCZBcW9jmejegvLBbeb0AyyeLY0RbyVyJ/ibHrshJb1l3M+ZUF
/7BUdXGdYqsSm2Iwg61S0Weic/7yePmFUjo0Lphy+8bkOqaw0cJAKR4RMG3kaZCJzTE2BmV04fL0
bussKhrRs68567z8HLGeZbJcyJJEimxD30kSzHCfiP2P70epfjjPHRIp6tWOiV31ZhSuGkguVApZ
u7sLrQT4/8AREkwmqT4YNOBcIVt6uditTKbdXJSl7/Z/LjuPpvFi17s2z84QpF1rbPc9L5VodbQ5
2k8Ubz9ngz76JMTnUFCfK5pAWL8s5rrPRI8sUwPadod47tN4rv0agiv3sArwwmBRrJ3a1LpaF+Lz
DgUSnmBrtRsz/EzeNuerWCAUBStkHdhQjgAhrI8FafByU7quyyijnRzJidcGJy3UA4Np3+jalmMy
gVDED8X4hAwf8RXHlynT9ZOPz5FRPoYPz0vCxfFuMOVcyDL+msEd96FoWpDKfKEXg+7NiV1ALtSf
GiO764azCbuc1Sqtws2bxrNHvZX0If9stJSbYpCemt5IbrsroZei0iC54fPNTAXjGn3neGDQC5pE
7kLsATITimpJ5KLD3SWMCmo6FKTCdrhCGTFJVpfFyFHRfc4sfdEzrrLIzFXvcCQMYz+nqGmqC6DQ
22+5VbItA4ICy9os758DnHqMvaEnP8wKDj4nKejtkdRjCuuaZ3GOHCMFBAarAL1NRJiUSxEBu+6/
yUgz8X74NADXlnL30HJur6juxyAX/E/fc0ouDpxADeyS11cjyfV9ThAq563iNguyWXd9fx0B8kxw
07h7OdpT0jVHpnUy+0YDUoWIsG509VkBmSSkQ3Kw55BmvxqkfvCj5CVbalTM4N8vE8+DZX/yvrdB
S4e0eK1cu9gRcouo/ObZ6jlwqv6FLQcYHdjAOpJ/QZ9pk+Knq97EgTYuaF6AdcLSa3PGHSHoypZA
ybyynS7KiC/wlAckfVrGs0KCpVG+Li2bcjqRyYRGZ/pqyJJcfVIemvSRRZkMKQb6SgY7PM+aHFGU
87JsG44TRkSei4iCUJVQ3FIFMWcRUPm+ZgKHFY7ez6srKmOnh7D4V+4isFsYgzUzrJA6YjN4qyRa
0FDAi+4RjOrCTjGoFGiigozqAMoQhAzukz/jIxRlPbfpnZpE1vFbwZnsLgQrA9lT99WCUvsr/qZ0
rtDasPrakAUyJMSdTGhcplMPwHrMmRgSjGWx5zAhPiZf0Jl2dFK+OZa9pfttu8F7FEfk9cx1T2e4
q1DADO3EWNSsiGNkePL1Xdrj+8l6MrQeEhvTzrrIkosVf25SRxBeTE2tDlboYA1aUSekAXZADruE
7vOXTaFB0E2YPs7RoBg47HP2hsX8GtQQxrAkb2CP1acEOyd+HrCvHvrNtOLyXDFrnqnjQgAu5vS2
50d4dSfshZ85YVAzK5lkA9E8GRoytS4Y/SEMoMM7t1nxHvFqKG7NBvF/EkXXJnTXWCjvwRxNCerf
rfAr661fZGOVK5Bj/y3a3vXDiGOrGqxi6/h5MueULx31MW6d9ujK8aM+EPc96i67HsxT0Njj3tmh
YJtSbblt8/5L2FD/TcoxtH+tgAHYtz+XJ933Dg0pfELSuizdALXjHOJMmyuaK5FdHgJ3F9TDg5SG
2PiPZ6mq61u663D1Y4UIoyOLTWm8WB6c7Gxa01DjhNQrGwhSVpehc634jwuj1nGwqAsIBhw5gEAq
ZEL71w0GBhPgjBoxosrxtLWoPN+yWgLWrH00CS2bywkEdZz3u6Zk2dbNRXU3I3A0uIDHYpj5+Ndr
duXawbgXi+ioQ3kly2mW0huE/JjV0vec9oxqa2GiN3CsSs0bq8eHJmNZNNlCAnur2WiKZpAwITsZ
zbl20DB8foZ93P1Dcb69K+vKf5j8dSeOLwgYCPEAYHhF1CQX+xdU9sajld3BbJ4eWxAcbTC5jkuf
RBQi/At4MADQXcLk5r84dbdrj0WFZGV8Xrs2YOq0FwGrAN6HJdCL6ueJj7krGBvZMUzf+W5flDat
t9/UC77EZ1a6UQYOppTlnkUwVVwoqyTTtp5m20pcMEUPnazxiyjVxe5ZVgcJRTh28VEdyIx6726g
PJbVdp6pnHbcgrDCCayFFIsdlLWyKhmn9NvaX2DEQjKrG60pIncO4s4H2ACtpj6LfVguUHeYGsR4
KvUGSxNzztengzQ732fEy3y1MQtOUn6g/mV0tHpeMdOoEUwZarKiWj/Ug/m9NRWNyOrNnR9FuX7j
UL3pZDQgnc1rVVhSPSOpYcf1hW3hd7NWVoYQauAwv8X0d/5ykoNvqDyplVyJV62fgXnQqY8Xfmz0
XJwvj/nnFy6niMhGLe4sEAgEu1e0HMUNK8APPiCm96o3K/ZUDmLcYLFSZ6Lm5TusZsUDh/Pd6EQb
/5T6RG4tJzajKbsZkNkm4b9vrc/z9mwmdN1Pp6v8QLBxwoVhAW+qIFZE7CSmiwL8m9flmJYEwnYM
WoPt87w9v0edP6k/Lx/RmJozJC3tZJAkWa/Ww/QEM4xNPtA71Jtbx+p0BESYUQ4LrumTANskQpPT
qg0QD8w1Ixg1z3LoLhOtK7w01FvH2d+6uL63D+TwmMCv063K/UPb0/00BdA9LZQwK62m4OlamnZt
Ns3rXq2teu4mqc69ywv8LujIYj9IyIbUrHpyxn+3HIms6ERVLfOeptgoFyvrNrMALXLdiUc1zK1X
D3j9MtBz4UqLTTMxBNI4zAuTkpMNHIjPS4NBymu8vC7MtfHBzL0oPJx6glqBO/KuUhRbANAVldZn
Rw/VpbA7+/yqTkdFIkZb2n+H5930p9qx6ZSDk7wHIh/i6/1Awo6xSCxgVFvkOTMXfI620n2cAwp/
nLbXoCeyTmvGBVbPym33A1w++dAhbTOblV7KDw++2BZb/Yk1s/0YfwOqy3Psv8gKsNNzcg8p2VH5
seVFfGd1X0sFwlWFi6mE/UoE8L+1IqmBZOTk7caDwXP3lCIdjvlT7UnfO/GNB+6ujTqr6l9+EwGc
KqXo6oloi9tv3hPueNeKpfjwzA70IKxjvW1YSq6Zgk9vKWFreHLG0g0Q83iCYiwYomGNpDqLmPye
KZpBfOkVIk9ol7A9i+vSTCfZRQCtnnydb7YYOZ1nxDSb+SpJIeLW+qEz/rI+yJqAZNjZgcuxZoAS
spbCaJl1CGuZ6RlRixJ7J3ntN2veC9jYAq2pJe5ohtkf4s4ZdsE54PivA0UNo8s0gWCXSg7Qexsm
ECIMfNNDZqagqjU/jCV9v89N+UriZzpMD0KPSwN0iIYWtT+ON/xV79YlPn1dprQQlqf4MaZOiRM1
5XH832IeClvPjmPPCB9Wom5ilQiHUCPIOrdMIBJVk9L7cz5GWLivVv9WN+JZZX1za0g+I809rBYI
TqVuekUwDOGxYlpQvpsfqeRoWKZbFMGfhPPwi1Rk/oOvLG/842oiYuYJtgJy7ko+8zoSOtRzbY/C
59PSO+mwajLfl9WrWUNfNZ3gyTPOIk6+kPdsnd4q1WP3x6UgPISVRfTpL39NlOi3AkxkgCDWGngR
qSkiG/tcjHWJBOyP+Sr5wnAV04Q3rWLONUAZl7pxY1UqgecCqXDHe4mKMwAJaW0gXVlOsmxlV7sD
L4OjcuXZJXwKG2zdNipuR2dKP99qbANsrsikNb+SsobOKHHa4+gwT22P2l9lS1Dm9XhXzAWShgXT
98rioMzGBxOnYQGy8zQN/iK6ZrgPWdAqdSC1zzj8CN9pUX4vbxx2zrpF4I6/XrZZwK6t/tqmtgIC
OoVFk0d19kjwNyOuG+kShwbJFb6TrlJnF4cHGmgwnqww7tRukznAn1b33GvU93Yw8ZtLpRLLRmmk
X4jNzx2XVgx1GcZHGuecNk28sE1vtZgYh+gmA4yBYw2pVcDuQVDFLETITz5CPEgCigPiYtBowBvq
KJDzMcdLtDAm2aJbu0Tu+YbaiaEPH7yk3JOzxrAgOwLH5oct7/ebdot5IR8FlxyLH0QNGJWQfdbp
NFnI+ZuJxGJ4XIknbUrFQC/hrGFSGJGLNA8guP2NMQ5iy02lmf89HwZSN1UiuKo63bnLDZUcaNGf
rJ0H/cpBFNM0ioEGKuKLp45mOm6yZRl7ZKtwlZThOn3wsesCj73O52D6Ub4B8HpxpKszhur7pNaa
RbrUrlSOsRb4BtqC3cPSOrbqOX2Ns9zOLKgmfbtz9NL/Qzs1wOe41V+2FcN9bAxWzby3suAj2wJ7
w7bgdAyUpU1rB9G0KENGi5heDc0k2nUoxuq08Cdzl17FKkJy98yjfy8LwSHRRQ+U0h/7ttG2F4bB
Nx2gBmPFwsiOEUTRrM1gjliKxpCaYnWVJb2gMEUKj3VrWiMc9ZEW6nh+AtfEelZo/NmbgpAQ3sFj
/thGE924BEmltrwG7ZZHUt6XBgHXfriixKnK6R0Wwk6nMqZMq17WbbrTPgpjS/8v8J5TvSQQz8T+
bgkObquDpegBXJCoJX3fPM/ah0kAULc5G1/tCmGtRLCqRQTbvrGLdA528Jxp3l209g90fjlO2Yhu
t082jKH+nQb/U3Spd46MC3N1p1r/smZgbftCcOU8I+hlbWtyxx0oF4/dmqUCL961wOyTbXWQow4b
WcXdBJnjPiq6WcbfYmkE1ypgABaJp+w4d6pbRm6aGDB2cYYJ2fc63NctlqPxyDGGDf42AjBES9mC
ddKySOjE/1Qz/JlD4TizYh766JYdxWwwYJ6JhKrg2VxnGRi9QDMWpqfTP9QehBqDKYazJy5pt9wz
q40wEEdiFDHvuQCo6CO9JBQCzbl4dJb5s+dwDbRMKr6lbwq1BeJIuBQ3kLNHMluHGRbmJsqK1E+2
Ohl04l1EtUFtleBjxN2fDwAQa/QewiCDSNosZE15LSiJncmzdUZ+yEIvWy0SCfWqnUfsKg85gUGy
gnCmYDRZNF8SZ5gTtjZi7/GNoepM8dTZfkffIG+MG5xYCCVa2RM/gKeWEYdOprJuqurS6jrkbE0M
QW/VPmyfpVuiEN/WHobS3ObfvOvmzapPU6HcJV9+p5zxOFvsIj1PMsMLJHqSSvJr424ee5A/Udn1
Fs0gUfnrh/XuPRt59TQX9hC2TB1Pnfm3G2AK1JIHutYJqxiJhnWNGBY77+jE4LUu+mMIpMrB+VzZ
5mU+77t1OPBiA0QhVkx6Gy9OZjUqf3dbk5TFtOr7TwJD1mlU8Cn7PZaMVkavxT176H2Vqrv7lT1Q
yLrBgPwCNhXM1usFrWhBMBKeIOCWb/1dyDZYOyODYvXJ7iG3OUM+elYBDjUyWuhqWK+Sc9YmBNqv
svyVJoJWcYlslAnD+KQEsC3t6bWZssKV55DH/3m/zb1Iyjky4woKY2tfyTAV24/VGlSH4zOYb3Q2
XWG/PmRYdIRM4BRmYFs4pPhXeX02ZLUbhgqtg5dYyNh91NMP397ASJsYeR7Mn50z2XxJgy2yunmM
++0cOzrQvSLpJSGzi4+gw/ZhRnPw/4oBLJ+KwXTBEcdM+Z4ny5ky1NZ4cydGJRz+lbKEpuXW6E1M
9DXbEyWT5RLdaSyasV2KXU/ga5XWcY8sw+/bPh0uTttkzfxXlrXMvL9Kch7Ap/F+WqpGqKrZKp8B
sJnhkQETYEZ45WCWgPF619F558oPkjE3Ea9b1zOFEOux3vGsCbnZBZcNBWVfCuz1+K4XNzOPYI1M
JjRYUFFz6BYOY4RHlKQKlnlXcKFKX6a89P/66X/qwjddvfp2LV0FhGOdIS08tKuBsUIl6JjZH1Mb
gSa1vpuzu2aMNLC6xEva14k8i1Mxxx6oAAMj+JdW2DR7dgObguYEhK2SwS9U9lcWqyK8KDFGRoNu
ti9gVS9deK1DwotxGOO7iM1wj4TRHxcFVu8iFTIMTC2uDqvinmcrwmCkUaDWW64vLMXWNeBbOgiS
silDHoK/0Y/eLTCfv3KcTonoGTcRRZX0VfhypC7eghjl/DieWbdf45BoMsG3BJheSGvuXuaDxpHx
sxbKclIZk2IUjWsI+N07G502nfXuREpiyTXvxuUNIOB0HTKfumgYZGIiJaAMGoAGeEqqL4KrEHFE
jQygu25McxMvr6EECarbOIGShrAH6INUJ3w2l+qwgJ0lW9GcdfeD9kSFRpmriRqUIyLrMjBDSS1I
+gVEPpCXAUu2FjXZU0kd1vFBqplUNvUlsIafLukx80tiRwKP5wBx427NxZgKBCj07g2tK7x40veW
5fkRnr12rfhkV/PxQkHGs3ae1bavneBnxr6y0u2Wb1MJMwmjPrr27gMkehOZRTJyq3pWKVcgFSh0
6+2p5GHyRwoDVLBlshDWCF3dttBWQBUsMaQAZ601/vsacjY6UclCMao8LpjS+aImGHLKt5nqlzQa
vp7nLuv7y0DfE37TnPZ2ofMpRdfG0oaxTQ/DOl2hxoQWxvLbTt3FGJ+hSvJ9fXDh5CuyuR5I2Trw
clt8tgYoIwYqTCfTLbU8icG/n4X2M8dHEwt7nnyUo3rZWM4CXAkqA+7DnqAB0x28jzVvvP45ojPq
IsB9QBcGvCqyoFSdzyAppzjFTc57VQO/U1/ZrB9KkGfsjFwrrJ/lJcIsxWm4qXMP0Y/7GBBQBdR3
rKTRZ1XNHqJh0dhHOnt271D/tXv/X9ZL+r2EQSAxSiaM2r032+vE9DdgD5YZVZ5ercY0lWPje/MG
VVaPar0zCA4FxHvuKysuU2l0pH6SMfQzwktN0LjcMmCLIpp8CRQoWqUopuW9t7VUWiBTv6w2R9ai
GNNlR0FrYE6Kc0uM2nwdTiegz0kMNpFGMEA0rOIiYhPb0nPBYkKcSoTHr/o6xUOrCS13jd3lU/tG
D/qbnxajhKajM0dP4ZKhbTaBrvbVVWw4inLUoQUlthreys6a2lt4SRAk8RWAO+1geX6MJPjKB717
hJztG1dg0slv0hi4Fuxzzc/NvUwyxmYs3/BxfFb71noYdjvdYXtckKu62yOyE0SUAFIjBaXT2YlU
Ayr5vBp7pmIFKeYg1DVS8r9+orP0rA9DT06e3wqNLpI4zxIPAsufKUvCb5ejX9GiyiqrJH1ndKzO
BNnb8eLiyKk1gQr6MYSXst0mps/Y2M1PojpAY4kSFSWiPDTE8B+DJDjoasVeRsmNlZ5svrhqOUQW
vJutZDVcr//9f9Lv4ICUIpovP15VaT/LNS/iSAPtOJM5jJQntBfEiTGif8HX6ycLMKKxrgTXOcBD
zTUnQCnaOCGQLMQHQHJCZ6L1RYLmFGiTIXBxFGhhmy6o816DyynpUy/bzcxVRk1kNu9G+0k+9g0u
5M6/73sTyB4NAVYF2x3skc5be3KnxnF9yiutiFaZ4wWdV3t34+0D1vL1Kq0Qa5pAB6ehx9lPBTfA
ZX9W3PbQEAxMOu2dCbQPKCogof6rFq4/nCgj1b/UY1hHiQgKpdLp3zIvGBmHI41kpxgIg1slKvyS
85F0v1WKCVXt0idVMXya4KWEW5c3s/ZnwPW6y9jgtPa0ctvOgjkblTvIHz0fpPC9PuaBmV60ZZm+
lUCOPnHpAAT6pdZ8HLKtHY5V2uUeZ5RBzZSjc2YRjc6LI0V1Y0j/G2MkExUO3LuQGlkz71+eja6l
RWS9lRbRe+g9DoEXvb3qhzTx7Hvo8tmCa3NiX8f/Bzl5xFpGbR4317R4xpF2ePZHLA1dwxYfUHG1
fdXpQDc2BDTLppLEuCD+v1yg0dAKJJwObjM68rfF337s4HdA3ynNH6QHB/tdJRYSWzAqZPXHDfrz
hCnNbarnbefmi0RJeZHWZCzSidlP7iEmOB01JpVL7vbqlaTe89mtOwmbny3FU27l6EhWj0Nc63tu
9xTINfPJypoWpSsL4wmCV0tgDcH83CAlJVhc7s6URgHtDpbjtTsh6GWxSb2f4KmzcjumQjZxsnhM
dt+7U02FfjAVDgjG23Vde0XnJozb3IaAXez5iINXyVOMIOSxuv+93tELs4dcJNEu3PzMLj0MWL9Z
c8aFBa7u3p/krtiiYN68odB8zdjBOJUQ0ufzv4WTlG712uIfP7OvVtEILpdK5sT7SQNuDMSXhGA1
I46lWx3pid34ydiKiTIH77PlthYk3KKL6YFHrZt7BxO5MuX81qEQrsekMTmWj9uEIdSbNp8GdmKX
80WnuVflTgEfJTmQ9O7XETejzEDC/jGMnx3kYR8Hh+oCzG0E2aKHSyNZ64M0aCOAhJi442qmbWqc
NcRIW4tRpKoaPrVc0ZXnHlSBNmsjnMhyKA+WlrM7kgpux5kj/1lzsAw4WPnWo3KYvtjimt0Akm6l
cuG1RsyXgtlAaWUu2Ic6rN3m/3MKImESHI3RUBJPksp9rLydLnjhrrIwwONUY3LnVZ6l95u/IZuB
/iIxga9iscj7oXXmM4Y+/4cKnHJOq6GzNfOVKXvigxpvfHNKWAP01aSUeH7oVCNJnt5NoWN1QO9j
z7O28Fkr78oodjMpnimUV1/LWoaDYFrP3oKlPMQ+ONvYTPFy3vZ8GXrYytHf6Mt1WSmGXgcESZSn
U+UcCj5DiM13OcblqX0kC50gV9UXN3a+Ja7B1OKrdUfB1zYrabYZ/cYHYVWxfCnmtLrXhynQP5oM
2mzRxMz42SUaduDVPQneUJC42jbR0AbevA7ybDSauUiqPFtAXxljmTmzGbhs0AJR4kdT6qCPAAsR
zt9l2KppDRL7l4Qn4mUqN6XOdY/plTJ3yzr+4bwsGDOjaCOrdhYsEMcH/Cypqchihku5B0vDIze7
XfQ7CGIUR9EHPz/O3VvO4ImwRhR9WHvLM2RbCiUhY5/h3PBdSKnkobXN5K3Mt91lfcQV4mE+zjZC
EZSOSXXqN5hbWYPBMKugfvsKLxh78LN1ILawSLfVx843kuxORPyrbzAiuFQ4C7PCNrlS1fvUqElN
MjRrR4Rr98i4ElRFb1cAUNqI9eqzaHfBhV3hVrcSbh/dwrHnShojnZhw2M2dKs1UZobJObfugudS
p5CbgMxmH73XzKMb+oSvCeKH8ya77ofG8TfdSdn0jkHg4H9Nja7dpxbcvd9VTZBaGmrXdFL2yn2T
0jxoQxjze7c2YscLBSw9h6Ma1EKbdPrJlUBGPArAVE/OHB0HYxZTtlTozOrsywwY0b9PoEy8Jtl9
K75k19SiM5Us9Uk3jsfAjAk1RCmNoiQHjJlklhZNvsbqJwIzcsm5HOpumVNHpQE+sfuq03S1eM3p
sdrgfF1PwoFi/dvKqvAaZZiHxx6OtPvXh2CNuZrpuhUewGRKr9GCZBiSdX100N8iceSgKUI2TTjF
KD6Ue3kBxiqFcZ5EV3ndt0UbLWAVkG6c6ans1Fuolz9LOYSZ9R+I2LLlht9IzBRw9+tV1y/mQ8jO
W+ltp1/RhDvvjUwXsODk2ZJROkInv0nXwF+Tkz06lJSt9QXSlkfQuHYZVPBRt+7oPNs1Etm3Lyzm
GGivnYoI6FFpu8Qa1P1FHll/NthfSyg3/7x7zIS8xliQi+Ov+JQt+dik+71A5sztlYCYP6uHV9mp
Qj5rxXUMg2xn2aYoDdFG5zFvde59oxMPbTpFCVFCFwaixeTvFX8u89hGjcPe2OZCjCTANTs1ZGSG
LQgIuzYEe31efcxqwBeue75SFKOp45LzbmA74IrlMxFlJY5jy+lgSKMNwp1wC6JbikLXVRCqfK/V
v8Rw1TuzdKvXKI727tQd/hHPhruy0Vy1MsbPodpfoqbRhFA/w3GhBaKN17DWqHvK+kB/w2jwJZQX
mxkSfPGPNFW350EAWEO/FgHgQkHiKVdcQ1ElkpuQxH5Ow3wthrWv7XgPTEe61Mt7Dyg0jiZJBysn
Z7cwusK94cK8IKYrPdn7NWWS3ls4d30smuVrGp6bWMJLWdxKELpAtvRYQbULfLvqZ8dubBCVQjxN
0/yW2Ulh3M7N3MDB7wTME0trWquSa0fXX9ta+OFfFeiD+PbT6PAibR0pInT6/vyyr5aJX/IVPTIb
NDr2uo7gHOxo4hIhkmiATbVKyQsV6agM1ODFyqkklp3ffxnojPCaoP8XWx0vKSq56DpvdiI3CMZN
M38WmXOS7+/1nK9KE/QustVjmRRuLlncL3cCTnq+tz19xLK+5oYyUDMfewFseR1EHU1AqjYbs516
fFQ391pSK4rBap8Wu7BREPo+ZtuHtUlKh5vzww33tUmusW86G//y7ZAU3ksOXzuCCE2WPd2S4e86
AILORKcX2t+jjL14V++on8wVlgo28wTqQn+piu31t3YdoSpP8foT9woeVC9ca66yJWkQCvzi0EKK
87oCJHRa6oCkNkt/PSMIRw4UeAWUnxlwQ+3OgcqGB0CmZcjTbg/7kvoZPHznMsLBA2K8exFRqUlQ
YSz8IioooBwAUlXZW2wKJBpk9KaUVm2FbeKRC9olLmdc71MX9w9Zbrt84LTOtFydigGcOPqI4g2C
YndgNaTiSEaKXDxU4gjjS78Ca/xrAEF5TSci4vWdrycTe+NmfNbNof2vi5qFZwsW0zdyequn/IYy
jlP8X+uURqo/lz6dbvdg2vJ8bulCq3eRKYb3Jvv9omiHl3s1IMt0Vzz+iaKr4Mbn9OEVaCMlGnek
aV1ZxSH9SUUhfwHx9578PUHVoEkrhjiZqi0sW+S42qBKKwuQHMZ+VsybOTOYN3TSg2Ioqmx5yhXo
pEhyeiIFvRHltbVpQRPscWSO0DZEug+yQXMXS7gthQ3VgCMcff7vGtd9zzlNPLV2ntcfhElpm+Kx
1vwojd9ckUyzyvZ4Ofn+AZmYWV2C19h7w89vsdosAwAJJXOnascmc0QEjsEvyeHkKeHYe7YAYo+d
YjQg7HRkzwl6IGNBU4+cRjhfhUfBB8zqaulqdlGNs/yM/kJuPFFzghsGX8ijoVMlqlzSHZvZ9+LW
Pq1GVPJscC0Kazg1LXcHvvMUxS35CKZr6GpeZwcieB80VGUf+fxyxPvqE+a9urYG6o2PuuEr4cJs
HRIcZsYfVed5eQEqPNMwJzwnUZnNKV0BTlO7WuSi4FTkFn+G+tP84PVAeX+M1N7lVZ9/AieUvPcs
Hf7WY3i1q+sfnRqlETQkodMjqd1POWJ8XudCq7R4+uquZ3NeN6Mfg+r3APYOsHtxKN+9/c2QWnyP
1qbliLMPcgbAKm0cDZ82yS39pfKSOTWdSjAxJkV3YCVeUaTPbQ8Deu/xKsYoXFEkRjkG+pVRTUfj
rpFnX05yyqVuKjW9FqCAF2I6tylzVE8onHgDAxLUK4AE3kSubVikvWxghm7DUSfuwaaSwaBgY6Dk
2ZP98P9EFBkORh96Nds/bPRL7uveTQ0149TY+HABBByk14RcJxS46hxwQN73wEdwPYxxCI/wF/+O
LU4mMhWGLE+s4o4RyPyovfoxOulWJlFm5kb3QE+gG4RswjcJ+i/5wW5qbJqkCwny3rT8xLf/1i0b
uYu7VuBkQL71A8bnzwRankePGxjZz2/rOhCwp9b0AldNGnpSqcH89CYHCEqpkOtWOscA54JuaPDI
V+KGTcfiRv/ObOLMeTN+tNcRHdn+yYwZOu+sIoPZL4N9kdguAiT113MqObK1LznCy7ePXM46/e6c
+1KvmDJxTmTg+G8qKQxPFFhJWOthAZIbCAoWRa/DCJaQoeeVQ/Xnr/94kfjisb+0QIQGYg2erjjA
p52Q570SToVnhTvVuHn0geC23rEt/PwUoWcpf3unmcRBZ1xs29iDnDFEkaG0wLjY2CnvCcqPgULH
1uoeO9OMWznDAqN2wEXKu9p4si1kMFgxBEHtjXxp3kSJRBULW7YDvgT8tNzz1IytERO3kjcxgnC9
VzSHi8CaVUiUP2E/W72FNcqm+7RN4G1/7E/qVh98hYAw5FHZjUUYWnxSa+9Lg04Zv2LvpUmH6kbE
oM65vfYXKA1NgzylXGMsB4cwP+XMYdQYtXzNmCt4yfN34ZO20WXoGgHJJjg+SPDq3mWDNZSwjVk4
HfzZTQuUaLdHpFijhttN+c0BYuq1U+/LAGynyxoFNpbJie8FE2dvu/HMwFuvy4we6BtY/Cb4rPja
KDeF0R9Mp0lDtzV015iThMg0cP97PvG6onCLHTLT7gYiWwAuRUBllL8dDPEVRPHqqUGnPEysdXCM
mLX7q+x7R2MuC8dL2Bw0Ov+kyzGdtwF8eKifV48PnkoyV4Vxglci6yFvYm/mPcQEtfg48R7h+NH2
vU8XJaJdMOw3+nbjxYg+a6G2wsvHcTLQHm+WKPG5o6gveQmkVG9qGwfJublQ/oLXpWMoKlI4Cn/g
RznNy9ZvyG79flZDctSyHHtR8WSJo809R/ya6zJTzeyywj8OKHwxd2GChG8FcKxdlKecJRaQDZgb
NcQfuDkPAbFwKjscPEQwnLTQhrvr2THaOmSFMfAIdf470gb1FF9H+apA756NfPdFlAXlHvDyDQtX
tVCoPTagaIeJijJNYveDajb1bQBqxhGyRmMKvDdRj/lc1NKagYEy7FvhRrB3Md6pLB303bFrR0eV
pE+79+IIRsn5jWWaGID8V7/ZytQaNtr5xGjGaPBTF3h9FMc3Uo6fqvyhp4d1ZPlRVf/FOmihEHMW
bljDpvJiz2fORG4JGEW3LLvAVeaN5JUnyvXaN27J7YuwT+N5nf8uUQcqpyajBb9QTKyPdoFC3zC6
hAQCgXqv40s1s0R1EYitHn0NRldtMRAiQOByTWbD5l79wXGofGvQCINNiKg9MWzc9eONr1tTONDO
l6tSUWUATVYTX4PmCOGI4O6YnkBgBzzwjM4XdnJVv4SFKGASPvp0VsrW0hgN0fvhFxenCrmnL2c/
NFS/638GX2EumHNgnSg+x+ZxGJu6o9iWHScv++qd9HhROqBFTXzHx/oTNJDfhovWCv/BDE5DHLGL
RVEnunsu44ESRtAjdGVwm9Y0Uslk1E91pdefYC+0aaf+QZDXnhPbqyDH6H1kJ+Jh9gfcyEWaSUEu
UUl6AdMSMTg66zCgS6NYZlpWP+wbAr3oIxZZCaCd+G6xoCVgn1AooF6+akCOzy2QWHa0EKKlFHE+
A65jTdUereNMNcf+hmkF5lM8CuNlJaDEDWUVv847/NGW9VOXa8fFG9d/G7uMPz41R0P5cQX4IF5B
Iihl91kYrzEW6JAsf5Ntr9f0sbZ+x4WfHCPygnD2Dd6DAvuLOnuka+8OTF1bNjyjkMGRQVhO1mzi
u/sQV0KFaTp7FsrSY9AhUXWw042FxeoPyfPi0BoM8h5YA2pKuEhbaXb1fCIJhIMJk7QphqWJsGQt
DUj0BNnRcsVy6FW8/hFnsj4L5AyrbNvWLIbmIb6sTCX3u62Sj6zbmid8hp0sQmpCB6BPRA7+DtZ4
eNYTyF3nP93c6yQMx/WT5xRbpczTKlpjIk+YHu4DmlHn5llivEmG0b3aR8VLopZd7BxGJStmMqGv
nyM62nC+M4fYp4iiS3azlc7vUJLmxyexSpNZTblawBX2OvkcDtRlCT5MloSEroWtDHE/paIncub9
bxntuURsfzZxR8A7QWatwV4S1LAvReFuJpZNLEKBGXTLNTrZwdVugQLZdA5DVfGLZnYHztvGyL95
+9iJeD0LZh3HCZeq+uzqkWsEeoSE7sS4Bv02bKk54uevSqs0KdZVkhw4fHSkG5TqGZLDrmlXlUK5
IuVe4iFL+VdXIlZPNNmF/Ap30mNd0Xjzbyhc4FPK11MNSspXuSwVs0eCv4j7I8vAE/o+TcmT7i/2
grte/jxZ2ph+i1QVxv45rkf5XBxLFPj6RKUlbLigwvJXQQQ7dLPztIpnitNxb1rqa0LjpWZ54re9
oj4CslEnAm19Ultxow9jQhPupBY8C0b5f7CrydW55F16G+dKGYNYvPNMt9KKxDfiJeHmZvHx9njn
1tYQIzGWhk8UnR9B64QuyFHAG9eRqnKyhMH2kCPu7yyafGImhP0tOetkKhNKI5U8YLoiKuQbarYX
IdOnmMi0ct98wkVfcIYMmLXB3m3k8f+HfctMfQb12Y/b4YOG7U47805GsvEa/KJWrWlPsZS+Dyho
ev1WEPK65QBwtjiSKJ/fs4xup7106bg5fT/CROx03T2zoXS38/rBKMAF+EABvaHPYVvdrwd9O59b
Msk7sTn61iwPhKozXbvXJWsmYapFwlfX+hjRK0QNfLx+NEqFt/vUPcoRysCRDYbLjYQLOpTelSIx
6Lv9SIv4l+kTCm022aaFeSes+NcrVQ+xHjIp38h7Kk5rjYRmIyx7hy2m93xDDHq3tikzuEm4AtD+
K7K3xkno97x+hBoRj9+k0ivTG4zsqwvCUh+DMKIB4hcodRWqi4pusjAF1ptbtvE8WA2Oqi09+sSI
wsjOiVHl89ueViLn9HCsvcyPVUckhFBgPZ76NLTmHuXp2OLIc9rT8lQJIMOWN26xXj8QcJoawQEt
64XZFnbfM1MNRF3nUmTcIhrxwyRfCxKUR8ipfvjg8zFTL1q2nwWgP4CIAsVzcq0PYysYDQ+O2mA4
+dM9qC9Jhof1nBbr+lDBWCp3HdyWrfpFek4Q6l67v1w9e9RbqoqGazJRVsXxzllPyDnBh83jIS80
lPwN2PWu5xdO/ByDhtDDyteYDHq6Lu3yCMYO8uye5xdGvsPyixemE0ukkpRRHE7Cc1MFzcyKyBNm
cu/gVRbR+8+zxY/iU4je6MwRuXVdYJINJKRpDaqtnXHq6VbbG6RXBjMvmAyFdiHIOqy4VrqxKKy9
z3xPPcLvwPAaL3fKhf7HGCuSHZLs1GYmAWaXih7j4GS1KHS65tw61EH0QHh9mvaSjlQ96it9/cst
vHyn3xAxFshcNkCkxXC/z1IyQ4foJQOfoaz7XgID00c08YJcddhEsDENqlEwuqBRTC8OiaCPVVl0
83QTVEDCD2kBipHkZoSwSumqE/PD+bDzxDSIQP8DpH5FTfDG5TwFdCi+k70xwn1fH3KKfc68Mb04
i2G/NzQTVGrfPIUs8gYd45szm2SlSrOFuKYyDJGiC0TbAGI7KyfJdRE+Bb48b/0NWRw9C9AfA2q0
jvl3CN8VwI+3jP7ETJUwuyMmm+43knBijCnbaE7KvM54eq3a/jt2EO2KIW1uteiEEI2iSWJp9O6Z
pTh6s16LvH6lXsGi9bIqrZIN/eCSj3qbDcu3reCRgK6uYOkVfdJLVE+jsOREg0aMCr0p/oiaVY7d
TbuIZDbHKN6gfes4ckTHI6dn/3q/np6w09FVquNtWfWbItsr2VobnPrDcfHbBk4nCs814EejzHs/
as2jQu35JfYcfW89T+dbPnZCJySwdif/X9cJGIUJFRvq8m5aQWETBDW1jOJMPvgL9CF9dFGxKpLV
NxVx3QXyfXiHLiJOULPnZ8wRlfOz6RT8wsPGSFEZ69bjyIcxBo+BZd4lM51luLSmoxX2dJVnI/ps
VOYyGNot/8doDYMLjP6JkCwOF2UlNSR7TaN3DyZnDjuJMINjxZMMnSlXvIon7MHlt3XDfMXo+Jtt
bsMMprLcFoegcztFCJvZNIIXT7DTQ0VGNMKDAcqAmwTId4SyucnLyxjBUnaqHQVHbChTKNV4o4/G
lXvufmiXtQh6scpk4aeDOJaYOU4djmKQOvTq/aG3WtKtCw4zgYXWAkAwvrBgiYt1/fnfeufRb3bU
Z1SDyMVxAqE9TY94p/a6a6iFAwXVieVA+Twy4GnC/UQQGH8fDxNTb3nnmGOgNGYTrvUvSj4P+RFb
Z96SYSljWVyNW3j4gYYinGdYfhW9kfuE8I5x954tM1vneHW5LN81JO4vlIB5Ia3VmEfESoz+R61/
yc8iSG13IvqmkBhP+Tr3X3YCogeaUhz48hh4cqzK+8TAC8IDCZwHJqDfW9zSx8/ue9BC0R+3V3kC
eKuSBkIHUV6ChmO5Q8nqYuLpvJdUaI0acYt3RixknYOND47DEqNZivhwYLuOMOv+nvY8HhgSS5DJ
08uMz8C+4KroSqcOpAkWjGOpcgyISFhHResh3V1RDbe5YYEv5suZhp3vfiKEUfXQgCVeheRqLrg8
ll1eq6YVV6j5Q6OmSzpD9WaIkOncQpzf/fVYh3joCjQtTUWDP6E032dz7tKXsbsMD/QCwEUR4YC8
UerMUouYYhprIxqVLKcXcGmHwG6JO9r7h5NV6ecA3ZY0pVkMpF4rgFvCDO166hIPu8H2PNvBrr/7
BaDWeC79/v68j6btovW+lbVirOXZOkbvrCk2x4GZXoKbRLllNDfOh15vfu3A6QCnYtelEUXZYFC9
tnxJ3bGAMDujvqbZCt29X2TIyzseTR1hV2+QLRbH3M4XhNwYiatvcw+GfnnvyxVzogHbdKkRMTcK
Wi5MOraqmFJQcBTW0LKjf0ISTTyptr/c2fLiR1WK8htQnHWiNv0YHPqDKBch0olbKsmNg4VR+yDM
Cqy6Yh9Z1JBkRBJ8ZtAFDN/n5mlb9/jsC86y+cyulMYq1fvPZmlfuOCjYJmC+X9WWsRHVvNmqw1R
AOxjO4nK5v+a3y2X29Qoe5gwamIOmzSl9ZpYwrFXeT82I8Ondb2xSQtk05RieN2KQsTNzQ+WQfxb
vtmmwc1ClOEVJxqY8m83NFji16FNwXCSqSXlKXhfjTxF329XYC7Dek9CXGQKo/WYeFJTujLzqZtO
IgXsRMsKExFt+i1KiZfXIVaWFKFeoXKIDJCjoEaPvAP68WJ1nJMj8nfyQ+XTL7m33mGTFyAKsOZW
ZFqAb/GhIUUrAnzuryyYht2eqV5Ao2hVEzzpf3nTVROrvLHblRiUstVQ57yNenvOskj9Po7d/qas
KWkOTyX5Ni7DHmX/vVI/UUJKOZ8+hafWYdEcnOxhmX2xlx1S6yu9S58gWoJQp6UiGzRWWJXIgaoj
3aJyfcL81BdzksxJldGvATW0py+EeAE2l1cimYVR7WMZkNc/KFZGo17xpMo1ByvmkfNJGZbGg4hk
KpViJ6rETKWZdHOXivhO+AlMAruAjtwnwqRPKvQ7YC16RBGHlSMrJ8oD5iGKUTarTvm/78RQTz2G
S9jdG0xx/yP6tWmMDB599lOu2hwXSZfplEpsMQXeW4MrHT3YN4zOkLDKIBFKbgC7MQU/ESrDU4ZL
vjmzcrGKHvSyj3gNlhgQYABmk3s7Uf+OMLSylBBjrSAlYY1/JCItdbN53zslALAnjtCkCHFCYur1
8uU4qVaAENMoFhRvJXqX6ryjMZidlcbWIJNfS+9t00WAZ+xEvxj/isMdSO8FqKJAuoeaqe0ebTf4
6jIWB6aj9f8xBDOMr42EaKmU6co2oLdepSseS7t4jAbz1Bw4msP9TCOE3ngL9YsL1gLBpVurn9Rm
xTbcnTHC+uMwwGjqVEvi1s/5keWnG+ROw5AALq680mclsVPmyKUV+8f1HN5EgYdtCz7pPGSvVJ/W
/3lIe8UipLJDRhg2728N5vwHdiJMSGkRv/Fk7qduIrhSXgUk4h4IYOtgDCwP6wqdkGgn1vjYoRJ1
vl3GxTh8/uqULwg3KNThFlzPqit18Mv/auqCKO4yZabnSxZcYgDHM/yY6/pCY94WfOKAyP6bNLYf
UO8NH0hgRqyiy+BGXfV4fjgtLk5dPp+TvWUWdWdN7O4XqQ2/cLWQVvN0isjK6xAdybcX8eFrKrrX
vqWZuXWTPzno5f18Bd38KxXjdrVWs6gw3c7vROPQfZARPnDD5wKknCTIPtVa5ZmyGOSxlP4J0CBH
nOuDRit2PxUZUwmyQ2XVCvR9x6agE2HaxYn8EjJe85IU1+qJMvdwtAxdnUCzAPfRMqTEYQhn/0BY
hrU2yuH2eKnMcDpx0zDHgShuzPwyn7wEOYVuwfkuwANNCUWKCQG076EC7gIDU6Pv0ayh4sQYKNgL
ZpPO1UHZ/A5yrneiJtw/jd01rLtOiosCHXXUPFEhPXMfbwAqrbvprRFxIWumr94AnKWQ3Hn4cbr8
pYZs5CenTEy3rGao8irDHfkBLGxl33jJbmMaBKdU9U+GD02Hmbl1okOPhv3B/mdKYNk9rj8Ocq7O
lIblNJxynOeyhei+YvGSHD0UvzNaEU966ABroovdu5oASxsmmowU5in64vNP+ZzWWV29setinh2x
8fIU3uzTHmtpJGRgwl96+aq24T3AmNugDrMuNxni55uveWPnc5Bxe3Upo4ircsjShHewDFEIqi+K
wEZdwlDMS8DGiJyc7kYB3fOJkY4LM8DmOSxhTeBqEMqA6B2CBVSSnRtuwS9A5BnNig/IPLFzQ8ag
xKOtKgPjJowmwr3SzWdqI5jdqZJy3BDXZZjlamNfj3hVYb1vla/Um2rz0e4N87gWN5fYCiqeik0N
4AW9/8igHjBE/vkCCXBBpPAcphMMTuc0i4T8/R1f6zjtgKRS1B9j+6C2VcBdNBZOea9q8MNW6ZIC
Xiac1d3tj1uxRtwe2puE7gTAgJNh6MgtDdQPatW7juh+L14z+fyW6GK+WqbDHNMb5L+MPjAB/wpM
cgJEoC+S9iNtfbzi77LDkRP5RoHvu2k/wPvZTas2lzzpQ3EFKFjlZH01CbKT0+RLk0r3KThLn+ZQ
OcheCpsAJ4EsHWH/jO23j18FrgwusaDJX2Hkjs8Z1QfxCRaaZgjrCXbjTzRVcgIdfGWzrmTBueJ1
y5o6+HyeYwBVWifuZWdM1R6AA9QC0sTHjzQTobPxtQpbyFotctn7bSdBpfFsZjdrcOQOPjDiglj9
u4Bgg9Mwc/G+vVEes4CmK+pYTfvW1YI7XGn4vI+KD0nkJpvQIbZTxfy5fZ0xwIZlcqb5HTeGuPp9
3ES2OmV0eWU4wgj268xv0fRxuphQnQ0AHQ2CB71esw/qyDdXVNRtyrfV1EcUC/A6fPVltgnH8pHk
30iW683U6h+L9ZDGcqImXxwyWW695w5B+r1BZ98IEuwtH7GK08wHY2sMsGP5b/LcuvUnCT8YQQch
SFpH0b8GOgcJKVVWjxPnqXPOaT6m3mUZsZgmehLTnjwD7JfY72VP+3C9buAvT0Qw+DofFgFSzjFv
DhmcxjzLO07aT790+Te+r/r9LxgPCY1NA6jGf1lWmXga33wo8ISStZRdgvm+b2GKozXyaLBTZZrd
Zq10SkgyaSFevpkDH/ZwnBgLbuY0YNYLHYBVGXT0SYcgt4jxYvqXPwLK0DhJElRZjHDF9YIPoOyC
Cg+LzcMowZBO3x6fSEfi5fcBezA8P447pOCShLgXewvFpHVb4MjYU2MiISrwzhdJUYATTm5btLT/
LDO8E/ZelyT3C4pi/4VAg2okzWDRdh9v3rdjUiu+MNN4KyAFfUpAibwIBmkcvDBegO1teRbDqD3j
QvceEaWhrTtlH7I4dJZukjET5Kc0MfS56u4oOA0xV+cEvFMluuBg6Y2Vo7Mnb1jJ8xgQGxLoThFT
2O8sykYrSxsj/meHKLCPlJiw06NxWwMpU/3UWFS4f/8jYrSSN6BNB82tH7ZxoSUJ65o/M6NpuWwR
f069NjyLjPiIBAgu10sfviKO1STzCpUUmTKBQLkHB/1moKGOmP2retzFCv1NBQ7eb1y0/2VIxR7+
WAJt003D32HQEzdqZVMPiw018XRm/RnSpuDnhERcH7K/5Rq6ZbZ5wjWbQLhqcjyyg10BdXTVddSb
04vMKa19mrxmvgCfr3M8x3Pr8Ph2bwIL9eM7zwCYJZxYwdJqODli26gKZ0Shy+gHdGvCPYgIaxn+
4dFNzPdCn6GR7sDtU9vWKvZSJsgQX2SNPT1PwGAWAn4D+TCfZ+jN6RmSTebAMJqhO/J9apG0kwug
zKGTeXamBP+67yzYMgkbJmsZSbyu6eKfKDu16dHJC4vh/mUcNzpndnjFmi/rUggXaQ6g9QrZCCO/
tBdc1wOyfCmKi5dO2G6HlylX7EfoqfxwRkeyxfCkPm4R9lDMbsgQkrP3Drk39rGX0Y1Y+U5+hSzI
7nbSevmTOPuamEmnDBBLgi1FVJz6T1baT5MQx6SQ1cJKRBRlmU9xDjk/oqOiNDILvh4mdjv8jFoc
noXTD4TtnFxEANCeVvbJl8AkGXzPydfe3Sr4Dn6GnHSD2OfcFsy+phOypSITQqlcuZeDuLLcWiUj
GJADW35k/0Oik4Uaq7DUpD9vQF0/4ET+cSfUcBczrzy9hRxjShSP4mXPypH9aUJs6tk4S+GPHzyH
iKGPhCNIPhh5XnnVdC9IgEIGkEXxTMxG3golk6XvgAWcigEkHFmXaPXkspzUSC5Yo5D2u2XGvgZe
dMKOliZwdaxzmh7JkO1JM/i3191AARCEmFkeUQTFpzRMmh6gsY1RnctMs7S1+Amtaxk78LrtwMjV
dodGNjLi8XdR6aL3jU0FfY9djhGLxsrJcvgnxKsvhFTgw5YFT1Ss5fXjmjUfjj4REqR5BJaAZBGN
cLlhURcglOzml2kWoqQEYWQDBhaXD72vvJuggI9f32+CSs29zrHKCEzVS+j19L98j0XnHXJ2jZG0
/JJLu1UC1lPtripXFYXZMDX9a5OoFS/bUgJYKFrt7k2FNsTuSEwIfktuA/pxLU3gndPyZ38Ac9st
9Bzc8pXLYaoQ5h9SHYAgiDZqYZay6aIOts9hVPBpP+SHNGL0DocvBWOMAYzQch/rawlZcroqPuMW
2CA54Fe+/eU6zVoMo3Wn+LfJyqQepJqo9zX2W+IbQKEtlZmetqGtN1EMPdtpptJdjFDEqHD68YTA
2MPFTYoE1Dqu0vHXH7QxeMlE5xgfwV30zexgSC5DgPRRys/EGo5QaXNx3Shp+egGoh0cWfWRNbR1
T8GTkDOM2c8h2BRnILAeEmUA68SeFSngK1pbiJifnoRKo4y2opCiPiYaHipkPn4DwjLmCZihlp/F
mW+oYmem7RH7BFBPlU6+yzaLV2lZBQZNhQDerARterKOQGK8nTf/MBFmOFz8yGuF5grSb3RT9ip8
z9KQqBFPukIVDGghbd3q8ckf5wz2K6ruRo2QI2capg8ZUYYSbIaSqyOQpGlWZvcvsqkWqaeVNpBq
54YGoLe5V5hfyT8LpgNdTyuIef+k8CVFb5PYOtFu02KvVWgRC8M++g08Szr1FDj/+J7CM8qN5TYo
7QR7HH2NZcpOdXbjf9mSeDJmQL/Vi6UoKNV3fEX6QjUFKEC1JrNcJWuMR55HBer74mSDLDlX9gJv
ZehLu2jeG4rUiIBpQJyji7uUWVkW7oNBoeFDpQ/KaQUj8YLvT94KScoi3AaOurecjkfEB+GnOPBM
qRiY2jWGENDjo0ctfBKFctLGOuxeBmq37O4PF6vQBeeAz2+/e/t4lUPhWyzlJAZ3uTKt8uvOO/ED
6Ggt6ReSQlp1jPTWdLspxKbY/ipY14PUMfaeBweQ+1ncy5W5bQh3hCgoxnkitlkXCkJXP5J+CKlw
4dnnEiaaupA/UsNIMavbo1wy3OyiLk1eAGaUgbbgLhJf0z7bYNsXttb5Z51+Oac+pxvVb+fSKll9
43n/q/P+G1OJBgszDeC12qWJd+faz0LYNapnXTkU5rRUMR8KUpFTuLShE/gtWEEpN7Obuhs4pb1U
Hg7IyJQQrKVMPBs6bLhcrXpAx9DVt4NdhNTOtc5yQJ1KVqp5fVpVIop3ELS+7eiG3vhx0DXql7yP
6YUJLdrCXT4kpGf6QPXP367kxCW9iGq2V3fVIWxBhvZjHbjQSWbOcrFfHtFhhEdbwcTF6Wr3LUR2
O4hBoznCwIc4hdMgaSyemOdE6TYYlFvxV6rt0G2LL27+Bbyg2TUzcu0LQX0X7DcPzDSRdQQrLCEy
JgFQizFMv95nK7LHcm+wRmqrtLBfP5RXWCJPHM5sB7bloH756j2K/v6o5gSo8PMYG3MVFR2p6Qid
cBf2XJ3f2sHyEWki7EfnIuejMUdXCWZVV5aOfSHmmMKQK5cmOkVnM/5FcBanA/iMbj15clPI+3cB
MxSItrdlryQYN1JzRMq6qPkPdf/w3BsRSVFByWo0pKaFxML8/J/9v4E1uSDuEOBj6dSmdBAdoMGr
AkmxNODmorlS3pXk50U0Tpsl/i5A5r9RRS3ZC7nGIUuDRGHyIVOPXZxnazoxo/5nzz6Vna1CfiiM
z5H2rSGJFP4ja6X8DR7p3sWRUyFqXoW+GrA14DTLlBvq7ANH6PiaICgixsFw+wG1YC+8Tya0CRGh
vBbzpyyjfIOPHG/fmEht+0s9qWr0IRME5l679+514RLcJ3SK3Z6Yxp3dqiwczDocGXTuw4bexl5X
04tl7XQNqI1z1lRHb9ceOSCkWVVVEWhoSPCOxbAg9TW+QvoJZTodRU/hdqObJ/1Lh//v0DczC090
44usyDV/PnaOSEo1tq1DNpJMPRKVoydlqmRQZnrVD2p8ZVWFk9UVw04hKVhXPAsTbKUl+rPFkCX8
4XALVBoLm50mKCfPPeJKoKHiL7XzGgfFnEn3SGFFmDQ0UKfpkOVOqH8p5gh7fy7gnSiEoSiIZvmq
m1GgfEejA0YIQA4Fw/dd0dGJjvnd5nXrw0v8pRI9GhWGDmkcZfN0AKvtS9SvopydprYuiIuJZ6ig
51JqYJenCn5gnNOw8hivsL5eqClJaU4OBsZpGgOASnbFracM3rIYqe6HxPe9sKmoiLIyFoV8RA9O
4+u3U6SL2wczV3lYTU1xDCa/byiTH7qkgmZqPFlTFCShH2OyLp2aXVJ1usDezEQLZ6EH7G7KBduL
hFu/7sD6QB+m22tAuuXaizzX+//MlmUaw7zOe8MfRUKptMYbGsZIcGLV5Lwe6FuTXVXSbEvM8jwD
4nufEUTtSZ0LtZFJiUVNnA/xGihSNKrW2SSHoDTqzyf5mPvDb2f3DbS6nPTstW7+DTjcGHVfPGSf
X/WrL3mCNkciFG7Q57iY3QkL83KaENuSRJ6vevC3vK/vmqroisGerfDDRzkhvHgtA74ozpoUhOa9
Ysf2C/HBHjap8WZ9ynw6wL2raGQ681aa4c/3xZWda44BgnIPGEJv5Z1SSF/wGWvI4KVY0Zcu4Til
TfCVCTqwYnoeCJJVVveKYeb9YgBHgXTVfaRJhlLeQucQnnWqDZzrA1UEqQSrFmMlFyq+pcV7C8Gp
d/hdYh3r+PupTjTyv6+nKHcFYL1H5NFofKWYB/aLEp3Q3B0Ks6XW/Caj7x3Njdi/UAfxf7aimCH9
ICGU2jK8/IUuh4fISCNG4E70Ms1811Koo7BayWZ4/wYyi3o7sGWIZBuuMq0h6uoCsl87n4LsoBSY
KUeTi9Nf/504Z2dAMsR6QOooZXNLwoVY2ejiufQ2b8jfdg1qN7zByEr5chvH8UuwCcJzwBNQ0wPP
Sz/CQQWj8Nc/QHX4VPjp6oBiU0Ho5T9JvJpJWURnnI3KaQEG09F7iRlaCKse8ROmRSd3RhSIPcOz
BheDATsSgp9kqpEASJ9WFEBwpn5PykD0mWvf9D3zv00AI5RS8nNAULKimA9Twdg4Flv4Cy7ocoj2
1wLBCIpCu39z/QyXp1U5pQuMO/9QBxe+ZaAuLeGjFD1kDdUsl+6E5nOMWIAZTa1ydEa8CVJ1EtXQ
ePdvanTgjmC0EuKMITk+0vlr6r0vbkUF0gsnnp0w3TxNKYOyHxdPNMoPgy3ULwTDR2JKm5WjrUVc
9a820R/ggtYweOW0kexANgcpZ2N27wTfmpBauhusjZ4fOTF/8YICpdW/N0Q2Xjkh+O3x+KtkV3bo
ZltulnWrKc3+8SuXlJsICwTSEdOXelfIY+lo1B+Z3Xcn/eeimuHk28Ylgt8zAkMXMmbQ7+/7hiY+
drmgBcgZ0wAqCN/Y2/ArF7/f+7pff3kIC7fOMwHG0Pd3Z3PqvugUXa5JFwm9ujgfu70Zkwc5SJj6
sqDbNuRmH2OrYg4gnoO8MiyFKXXYkaiTGxQmm3h41oSIaTbCIImclhoBTSGz+8vN9s53Lu79MTrq
5Jzp6EcM0iJ5J77ZfNG3nX3qWGgCwA4rm8ut5dTNDT7LOcT7pKyxbMk9I1k3LEahe2doglSBHWTv
9xgmnVW2rNJz0Jnicp57fMttGSj0rmkTZwBn79d+JjlIfCnMyAk9xdZaolo14ps3VubTAYRrBdJa
7jGZ9qYy/XQoEZ/PxwkstFUy17KRZ7sKm2YN6SMpyF7tq96COYtb9hxAxjkMPBLtcw4JfNkemaEU
xgGfm3KCNXydn8eaOObYdaQNmMxmQDftwwQy2lLaEf5RW2M6xfk8IbgAr2Gk+kVe42KGIqEYCodt
107lUCc4gX541ZEaozIIi4G+8cKTZd54K8ieWdyy9WmuEjrNOnCxbjd22vjYJOXKc0F0nKEwt1hf
4bnjoNWe1JhL66D7aEeat8YtTGhl9IJG/tI908o4vOHbloEc9h/Pqr8JAFDDYsw/a0FAnIjUnAWT
Ks29hzaK3qnYOhnuVFrdT7w+DzeHk/Ss+F/69QiSGpEhkwSN/jbenzZXL07FXVTYDzAwnGwJ31su
5sylGHx4qf3/Td1TafCvMQYjA+FpHdlV5LSQwQSyyp84NXFFaqiZKdXKRC27Gi4OCb1TzV8duXfp
0a8cOE2+GFRETlFpSuaZ6el8uOh11wy4adFFFWnYIyhvr4Xr++DIBQhW3lC7XBS4YOBrZTnYY1io
GFh+NYaCSn2arClI+ygrEmtSEwDOJ5aVUHlM+3hWStoXv2rzlt+enzMTgN278j9DBX77DTrWVQM9
eXl/gB1O2tzLfq8gQ79tumoaYTDTiXKrP2G/E2D0OqOPNrVmJLSP60jim3gGWFpZ8LI8XADKEdY/
25TQrRmanwitJ9VuNYQKmioRWzyJIr2qwv7gOWi7liAuPZt+JX6iZn0uitenDHkCauKY1jfFqWeb
dJ/pbzh28pyf15+QDJGV4lBFHqOMkEFqwpti9UE39vJ9RaDAW/WZAcj/Eh4hjR6m85zoV7os9a/E
fMHHxHObiVZb1yKc0/ASX7GaqMcBJ6elvSTepYM5C3iaIr8XsYtTZrXyoiN3ykTFXucTomk6yRLA
o5tE+epf2gh2FX4pqV3Sfa4PAgeWvs/QR5m/rvjUeDmPKnGE8zNtfOPbEYcTXQ5hmAC3iv1cb7nC
vkbTEJIke39/ZrVg4aGv++lvr2Kc9cRXiYWhCS3CBkNSOOJtRJojeGxzkZn0fIt1mk0s1CI3yquH
ygaUF2i4NT2M4gJTAuCP9ie1Je9Nb/FLOLe1VZ4lv0ae1HsbGdWBkRBG8vAsIk4CQnmNZr2fd4dm
3k22du7AfB13MFU23JcLlAPh5odGcsH6b6N40Tyc0I1XcnKOrQNP8dvkQ+xPEY/0FK6HQVDKNRib
XDYjFy/A4JH+Tkc8g+ykiM1Bbv6nbiI+AYrHeH63KENza68P97Lw6xJ1zWSj8HK1s68Sov/xQAn3
t4xNCzihnu6lRMPnKeaD7Xz2GpfqRQPR4v8tAxPuRcLOLS7vqxdhJqh3Su8RT3MIg/5PoEHaXEig
iWkfa1begwnY0W2LrPV85BUHdjY73FAB41TJzf8FAtxw3DVqG2CzW6MZepcdsGiiSP+xD8zQNg45
6odwNdlMH7PG4ZmQoOluzcVnpjrxmPfsOKc472sRnydAe+KeTwQAKRixZqi3p0WzeTRFnbgYbKX1
u0P9RAUlHjxWraBpETRWWF9IyIRsXiWGXxoLGRh6sWi9XOFQyO2reDLonqsfKQ6xGTAdCGf1xaab
B2lbxp/gWxAws2FzT1AcoRH+5E4fZ0g+/Ee8UnJ5zfZ5tsUQc1RqH89dAIQevcCaotCgHqBAJf6n
8ynL58VbUulumZsNEWHsAbeLVr/BRKc6M2RnLv3mvuTwoss4gE7W9CgrAQ27sxwEMX9lf2ffa4Ip
W0fcoKt7Vs4X664WdMiRmpCiH/sDDxlVD1N34qV2oO2sSYRlNaZQIbdvRjDC5K3jw42w19BYdcOR
oyLrUhkeEs6Y/4qJJLQDMuAWwQ7STjlIX32IipRU1avcJFyUacLrt7goe8T+lwcw4+IDoRYddB5J
p1hYVPNeFj4Eie9rk7PZFXr+Z/VYLNfVgEzWDRY0bmfoPMl0/cYdhnMz9wcMuGFHd2cx4cvG2Oyv
mYrw1vTpjFWDd3s3/B06i9dcYksoyBwdn2CYfzgGJO6eOVAL1SKVBwGfKwMC+dnbGd1Lw5nW0uvp
tFt2B1002M280du/PEiyc4VsuP6TyEx8w2cuuyX6FNA488SznfdefXsHRyB8XnTXzJK/nO/Q42zG
q+6KrIZpXvzCIal1/ePALY3lzp2q0YSGoLBbYoqRPMYvDZjpau57DLQVopZPLeR6UOHpeBl+UCjx
kGlaxnt2luzu9XSKpZguNDgwXcvu0zHUyUg9CgukG8jmgY99FdBZ09VZkQ1CsBKDJqKk3XZIjho0
ABjVGo/T10rdadJ84lq/JUB9q5uC51ElPc4MRUzGgT5KllztLGymqfWYpBdQ3dKaybxGO6R5vKWM
++kN5cmRpGB74SH7L0rIgj/8LTUl9nP5Y3UEYv44r3UkZ7UYUaA1RxRUlZr3KMbW1Tyr+5aZAvxi
LdzTqo4dj9/Hxn7AZGv43/Bg3RPQzoIMmY/4DGctlJxXmKmoyPTdWpL7AyvGsXUJd3ZhruenLGw2
NBJC53/KoAbXmPuzmiEyAZ72lqsQ96U7KKt7swa9qBKo+9M5SWguQDkeHUVmHSFwmQVkv3bj6vbQ
v9lelNjgM9r/kHkE4orFhFndimAMYKfqsBkQDtptNvLYiXbS0JatneK6a+jOmsccojo+FrM/glii
XE+a7teGULAQa+mFCbuq9IcHhjRkN2wpsLZtVUtYkifEdXHNn1cKjKPQpWPPOqpufIW1eUQ9yM4a
SGCeMbAiQzg2sOM1rygmulIH/zEK27n+V1R7ogWiK2Wa225xassxzJkr8/5De1N5XQisgtmTdT3c
Q4FiF5Nxald2mM2UIXR0YZHiSPcNB8SdnEFsua6AvCErRYv6J3eZA/ulLFhbBjYqmpUR2/mqJ9E2
biFD+seyqqlCsfa3L4i8MjvZbpAaOUKX+TSDYQJWbhKmiuU234FpXGnFYAmnv+z+q5pIighWTN0+
d/B5qYxxUU2Hc13X1zpdL5TLDJD2HOOK+sx5Z2tqHlaHYHXJGry9DcN26slYrZeIA/facpI3+ExI
zQJdkoBX4DJ7zDj1pErIaIV9lQHFmD3jIhnr08tgGBrgKu0T/BwU/YvMJpBS2W/H2vp6H+J8dir9
iL1DE/81BFC4ImvEnivi15+8jrNQHblGvQju98zJqoexpmXUZYTDy4N8J4PRd8TxdvDjYDAdApoT
gtTulf7X15thQlub5lfdRnV7zV036HaA7hpgnWLRXxuBPCrsb3zIS/ERBuZ24COxe8NFi+eyS86d
hLzqfCQlFgb5SeR2kv3mHURYnAnJF1wElnHxZPEkTvZLdmD8j/rYPuAP2gi9aWWO6Q/xfDc4Wr2S
SlbXxKt23KNM5pQBFvYz5Dnq+lb4aRFWekeS9Kh/3zS0oqN3uGgeoMrwoyJ9CbT4MKmHDtWjS/3l
9aPJw2fyhJeRNInwEQwQas7drtV3mmG8f4+dv54KiCMmDYcpk8+R8TrEOOIE2sJhC16vxXhBP5Ou
99F3y0P1n9GkVr6HRwho9QSWI+Atj0OW8Fi1Fpm0x//M6ZvDHbSe2lrUxPqxwuVhFZTPRD0E8Ng4
ENZflFqY/OmC99TRsHuJgAO5PnbYe1yR7NCuxoJl8WOywZ/0LE7Nsotc0pFRvf8LuuPeVVB1EWgk
FPfAaayy1i5BieCekpM0xkzLudzF8OM0gQGXdzEsv7XCAikdpD19hJFfbNAIcfdUzGhKZVFKG/sx
w91rtEH/UFykD8yP71tc7O2q9N9EKK5XGs8Lcww+eJqCZzNjRB6W8SvxbnQ4XeH/EvFJRm0Tu47m
B9WGtiLuQfGjx/9lezuh+iudCuLhLBs4YSfL+FihMAWPaFqTDiXM2XaSHFWOBvHDq4qWNqtCGCcn
AtrVyd1muhw1cGkKvBKgEZB8XQZw1A364PoOnWRLSHeqwvRPwSrafPMprCaHBlVyAUCLD6hPVtTU
+RacdYppJxBNcw82WaIzqy337Fp0jv/BZC4Tv1Hu2Y3hhr20xq72zqqxpUbEiN/EdsnOcS44qufr
Ur0uhxlGyr4O5az91wssTAf1QI7uDQIioLwglsFwyR34uh978GifaPz8b3Wa3AaeXlRtbYtA6vo0
Krid8YRJ1rLSu6jpfo3aVV2yJWQ8JDruuj1qYUqRbiCU4lXgHIP9pYuYg+8iCDwUwubnRYfPRw2g
Om96FqDk5Du/4laiAXTWHSsaXRHNJSU9ShaLFuk2gwe4jUml042iSbUtfBdnIzGR8pZHqDJvtoLE
Ikfg40WMCOW/ExMCCu5VoMivMx48IEb0dtU773TgKNf17Zj5HDQQwsq6vkNVwMrAbw9oDdcaL07c
2cVey19xkjuMqqrJyDbXbIG8oV7XRmsQnVw/YOvHVnEDHvW/SAPfCSv+n1K8LValZ9csGmbH2C+/
fs72zuXciH3rGAp4z7/4dkkWKQGrV/KMT+b2PKCV+QkmR08F/fBpfcRs6JshAdcqiiNg1oxoG5ze
mNdQB6Z7YGXZ4ccMDYX8c3ISOkkvo8HjPHhfvVW7FZ6hKLX4kFQ3frOEMKlKjwNMQQx9pA9rmkdk
27KOIeiJ7G2uJTKK8TGDALIrJb/ui3z1giOIvrkN5vuhSfOZmkkh63n/nYvaN3iDwYy07uFh5jpQ
ZSdshJb6NXGTMWODsgUEsYWBX5HgK+vIgyOQatv1OkOdcbHRM2c1UkVJPIUBigiNB0fx0WWRMx8j
zBTTqiCHPVJBF2uMV83wjkuePI/6MBBA6ToDl0yD3SvMB6zpiyM1oPtR0obX5p18NCWu0weuheLl
tYW4mc5d8AcyoDJKjltJzf4wHfY02tZC2FKBTzpblSm+WQb8HAJIkkhW42ywetuSvb/H78deGQAc
6m6QYIAwltXewiCwlG2okbV4hxT9jM8WOXonNBYY19vNEQiXDcGr9lHm1andimu0q6QKidS36h6C
anhBBXPWoP4DSyvRD38t2zJDfAUsBV2ffqDdprZU+GKvCrCz0c8QObgovPPiQazDebk6fOdf2QoK
nyEh+ke19snWslNhSA8OMuwEM+zE4eCe/x8n4ZXj5feD8wERNhpahEBEDgtWT9YgkP4qXTN8Db1X
JVQOGuGyMHpAZsxa+SctC9gbrYhMpDpFiPe+UrcbX1HqfIuNOkYXAI5cKRSgnb5qQWmshAlyE6tQ
NkzWOHdf/QTfezQVNc5Tjh05pKEgy2C73/clkFEYfKk+xL3K03Iz3a7qkF6BFMH6JBnLk0T8HhWA
lAvuOD1iqcn1UosS1LGRuTeblxCjPALkVF/9eosfXBSefVzbQzgCAFscOVpIYMOQcTlbZQC2Bn65
2548fXbcW+lSTFnxFJMFklvrFesB2YCAIxa97y9ObS5QwzuLqO18DWzduCcUzU6zXo1jWbUj+qxX
wMuiNgEJ9YfiwPCcTb2Bs8SCvEqjf/v8XR8Q5hhuzPFD/dA8Hvv/ADZYRMLUZm7zsQlnufXGDHjq
qCIx/pj/EgvIid+zJbDM3m9h00Ht5mgIbgZV3D24LC0fJAhtQK+FjgOU0a+avF5FoMzZE1olfnQb
DxO5ZfogSTKAENfJt1iDnwNME2v94CbpfPmCkKOdLFM1Tt0Aw2OPaGd2s7Bc3goBnO6LtR2DbZqo
ZaLeJ5zv7MPgiMbVf0s8HXjeyOiOYnpmGyZSXxThmsC9UwP6bURbJqEOY6tNc2ERpeQ2moY1lthM
T3zzWo5cAXm3hB+n3np8poWXB2XRJ42jKC8KPoKvyh9GBt2zcvL0Cf3YF5DGSX8BYRumE00443gE
3DQJHNf5ciiWg03VVZCRwFjy6H3BZfkGIg57Mf1s2/gic/jzry1tplem3QFoNsGcw9DDUNqyWxx3
hNCaSl1kqF8eFZq4QkHNFdmgnI1TPmNlchXb2OCC2uKbUtOoVRPcRGEoT2OH/5cYYo9cAyVD7xN2
okUnycM+yJHhYEF/06+9Pa7OaERmILnygevF/YiHozOCa4vCJG7teOgN9fuc8vSeQcA1DPjGG4HU
OOcDizkHykYdzMNBtvLsAH6LMRb2waSPOCKF557yeF8Qpp76cE8GqBmYBa/KZfU0G/aFupe0Zu5h
qgQdPYUPgwLbVe92xgZRSU7L2c75y5yaTBaCK+wFZT/lr0/9Xaxn437VtJ+GbT6/VYLnyCh3zjt1
acmo+sWru+a1wXLUElRw9ZnL9TBlr+IZpJY4RnDeoOmZKGpc/mEKeepEytomo3G6kx1D8wWLkGGw
HWXpvO8+arVnftl7pOarLcE1XqTAlKwyqvD1zogaeaXRPwuKxaWutIdLO8a4zg0Wez679UM1xuBm
8maH+ehW8JopiwAcg7jTsYk9CClruH3UDXA2YRx3gEv30uvvq1RGXzlGtph6L9e5zZwfaQpCtZCA
tJyPf/ex2flb8xaajkkZY5ptU2RZ8nq36tpvSAkZszmbYE+HxFR3p1P2/mPKLyaCbSi+JsVPoYMm
jW7q2cqDd1V3wGyVqE97L7+mwFN1vadIvOOkLWmTgBNgE4j5UH/UbRqrosDr7I0ZBcWdnUFvadxj
RHIRcIpiodp6VXS3Y7SxSUSCusxF+BQ3Ti6p5lvOMY3X/XsRqzUheuhbQlijW6is83xIQIlI+XOy
A5bQrdYto1QgnvP+O5mW0/lHLfMgqdlA2cTC+Qk9YxutMSHfRT3SoL8ok+CvlK3MRBTWoQQ74zsF
GBvOsyGN36xeajFIofgUPEkv3ZHSB8/WNbOQdQhE/8NHMygx4qqYPNVvL8jPWfKEmHRW/hUVG0Dd
hOrKETUxJ8TnRFl2whcnJ5SW1nWuig/VexJNHSncbdHgY+BLGAkhGq/6HV6XmRzJZa83USp/XVDR
gBOH1gWhwtqpxkywtWecwEIRaLky+F6Kypq1/wFxOnlVeMUPIQhciVnIilDmF5X5SwMorFiR9hSQ
pR5YXG7Jn2wSguKpXUp0RjoXeNbCuPWwt89fv023o3C7srxyTLxLvoO2z4CUMMgClAQJTI0rdTfH
GfhW9Stq5r5aTzozh9eYUseJID0Af5mvQb9Y+jZPTqMrNZQ/vHhCLRUwlBn1kZHTm4A/jHybtsGW
OPv2knaa/DvpHD6WtEJHlDj9kLOsWYPBOBVAkiB8oj4/gWGZgtYzI9DOm4JQqLi49RzvgUiVz6ei
AHYOtkjPEj3khk6QHECEn1YkCwFJX7dw0uy8sNtJChGVzcIo1eKA+GP4cDB8/LQh8zEar7hrEfPo
WKp7CIqaUFCqxfH3icwlmOy1+WTvs6qB+kbLKDT6gy/3wx7aucftuihUxuO7iB9ycx1KbK09eiok
0WVwcLg0ji/XxN44qvb6o9Sn1fr+zF3RFV54qCArvrcjTmPYsR2KRTv6kYIb5tR9uOfYb73c5/Rj
ndWuWgo07u+ajfujey6kQmn5tIwd+JYi/KZZptBufmCjZ+GdEWhLwKJDJKRbfVQOZNBnG5eN1vvn
DaHJ6YTxQmlfQSA3a+kC/296V6MBd7mjFbKmfIRw8YdjyRTtB9yu0+wBiw0dmHxgcAUGJejG2DfI
9SG/Ghbloq5fHV9PHz/B1xrboth/AYyM9T486X+gz8l8ip/6HGO8wJVQFbkRpeZchdE6oMWrnDIh
ZZLFYA6i7Z9oIg4oHXR9V805tBkroLydhC+3BWw4a4Uxi1sIe67+ZAw+wJM6egC0c7KH+VdGHiQo
tJwXCPGGzdKe87jFlsxzc3oK2+5bHGUbu8Hwp/c3EMjvaSSuHQXxciIEcGyOsptvQrsCB4PFEbSE
qJFhMhlDWu+efDrkFAxIYe7rFvuFhGg6d/TZFDlXqKwvyD8HyVLKcRJoCE92SS7zuUaA17wODDS9
eMf3bI1VNVeP3wrvEfhu6Cd9T3Bf2166Avp+CewsCDOmktd3sWsFEp/qruszJfrToJHt+bqRGY6L
+cWNQlbaUOATbKTsxOfSun/wD2B48GpHy9Foj8sE8v3mTV5Ez1zwPQ5HFGM7F/EoKmoxsfmknhJo
LkhI4Avg8tMlZhcemBZweJZwX1xFcUixyIDU+Rou3HbwjguC1ZH0U4jD2TN79FWVWyjgR7hEW3yi
NBE5JIYummY8EXTifvjlg1ZCCIL93tWHg4u3wmUuN1jn91Qu0co+IXuouNc4pWJhOmieJbjO/DvG
59ldxRwXsB8XODuUDFjw8EOgGQJoFWfnIW4Idnih2gKdINchoPe7PTwVWAGe8jrj/D/chAb7OI4D
a2OVOZFGSzouwKRNioYSmrf06Ymb90mu5E8C85bi0m3Mc+EkgTLggO8zWaMa9s5IZaIWlPcMPwtA
wqg/nEwT7cH0YZJ/7+N07WOFX+ZDeAQBMlbO58k0GHsERGGrblTE4RBl6aNo+moESc4hXXwlWT1Z
YIwGMMWRx5HT659jp+gsLkjX90td2bZCz4xTRVeIw5AMHQsppmWLY1qFcuXVVN7y3Yf0MDW1odJb
5ejDSx9+OYs6QoIwDCVPb+/W4YcwSQd5tt13mCpQg0bywgJtDbmHjPGdKgkL+ZANKWQzR4c1XPNA
E0aJLbu3SlWURM5X5ZtyQ87OwXjRJl+tqnnEcR+fLgPjEVBn9NyyWNAX1Cg7DWRrfS76fKHukO1L
dosp7nQm/HY7Z9xGYLBZMiOKSEDH2CmeR8HsoTiVU4PLUwFM2t/bDjhGjGcrytVxYRcUeJwO6oWa
ecl+xfslQluduwSRWn1IyaNvkwPZzOyNxGZpOfE1LpLLnIUc0msjlbBtUMqf2+v9xHRqXts0cowk
liyFqtjQWmTdeDZMDT3OjwXXj/qyxOueG8+95FscMSMOU5ojUe1Qv1lEmW2uBHV61mwxgUMWIdt4
txIpLhEu9kY1Puwzq9xMwFH4AMaCKkYxuh/SBGiaOf/htUKyCO1WMIVcB5xuN85DltpRoiZfeVKR
YIZV5zoS+KvTMogt9rvfej3SqnwU5o02nb2boGxFPPQl0AiIZ3WOyQ9m4AhnaCsJNjED6slO8ZCG
bvEOEPdO57WVM9Ry7Zo1UMATxUfJPNZl+ZojFgcHWvciQ77MlHfr9Lx6Hm44s633ZceFO22jaHEw
Xdv98gzUdg+3Uwytq+92pJGoCz7GVPXueBNAbW0iSyMxmdX8qDpfqiIR8FFqVVKZVvQWpXiEumkh
fWHLV+qhOMcJurpQ6+V2PB/I+oRHvfgIHrOUa4LlnUwBLNMMO+Ey0SstudOdQSVk06z628ZsPFeM
h0476FbMk6gVXeqvmqGm+X/PgtMs9y7cdgFmOXOUP7tVr/jqmXvEitfW+aIj4R3Wn+Iv8UFtGB9c
fl17Kb9jYDWaTKJwI4vY0dljHkBM/AMWDuUBJreV7jOxbWze01MouPEB11Q6zBtpGMOn6+SFJQhk
EhnnTWnMlrh28XJghSFCMKPr1k8IfmUKU+wZKHdQ5mNLsSsuWbVrK/ngfdhbojD2ZrEL5xvlPYAW
/7GlklHMXwajC46iFdEqg7XFFXySmpvYpc6Ruy42lKnJfVjf7/zpYFG41Pyj9crpnhdnA4InQmmE
8u97uosFGe4ECsq0E14lUpK2mpUs6qk21PHJKmWqUt4XRkHFSHa44pq5rylEwg9SqPETylwPY1rY
5XVg+MtVucj7uVlgStC+ijAZjRhn2VSz5bmgGzHRi57YtUZtets7vq7UJA8xAnu9lzVyh5bNiPxq
lu9ljYtE81y+/o0h8P5iRwz6qUCnJxBb7qoiy/L4VZ7NIiolngzXjyybePBuQBg03s4Ax8bfsFUd
tx6MojVOjJncqVpu+ohWfRKF2LHgHGqcjpqGWD0SrDMDZWepMk9Gwp0gxLuDChrUz+/g9TfMlmm4
ZiZwZA5isJsjZf4QOEUrg5BQcf8Lp1llM2vvmvtjB4v0k9uHMyz6prva+a1sy1CTbXHsShGsRC8r
WPME/AVfGPlhIF9KZroZLOWthrOFRENGqs1Cs1h+nmJQtv+ngp6PKcdiXlXxFu0BScbgaM0MFyIs
Q0XNyMC0DOCKDwNCIlurpG9cF9U68B69yroIHglQgf4tjmDvjLPWquwahXJPRgjzvUVTbdtoAAQD
SPRcT1BmAkarxo9CJx7FznSRegdc04B/Y7pDIOPmsEHbwXsNfUV8LNn9cJKh+3MgPLWe+kbylhoa
cdYYxqr+FuTEW3DGLGszIpMkHDRGO4m7FKE4ryUP4ZUWLdcanUjamVJWw1xV4oIawNrIG7A5NJUl
QUNdBSf4GeSne15Lwbwh7X0TRcGRx9HWqIzA1wOF6ia3vyYZihBnOTx98LK0Eh3h+ItgDCU/QdDr
muHl8v38lKJVeOk/iKS9uU/lzJmEqxZglhH6XvvFqR9KZihhad+0FN+A7bmDAIP0g6jGHhDctFzC
osPVO9awXERh65fgaADjIQy3yLHmR0vKh77FRgIo7wk/Ng/hCzIqkrsp5Uwve/l3DpnqkL40OOkz
rqHnRrNYG70IawzHdQcPIYedDy5rvCKPxBMEWG++GiNP8H48vADvUfr/QYbXuRjxefgfQ7QSh6GX
SHygkekEddL93IXyrpZkWluDn1hKZZiItbDLIV48bHk24BBlm5qfYF/iX235QgmPDlqqXmDl+prr
Vyu0bFXjKri9VbjSrghgdTPoBl7BUTxO4WE9IjzgU+u41oq8aNe1M5a/EoDCnQMU3fPfxSHRIQZe
0CK0o1KMPUxNcQFNfIREjn6ccTCUMx1atrrqdqgB7jBxN9LAbjeISG9c/yQbhbyWnGooeORRsqfF
v9J0/0u60iZbOcF16bUK/w4omE/ocBMl8qM4xTov/89Cu1aJNmcvHtj1mIxp45L931RkbDOHpcmL
rcqL2MD71M57+KOi9loDJ0fKsgrxQKnEkYwF2dAOChSFTrZf/ETPBdnYVKtmoPldATyr4fLJBfNO
9xYol0pOaBlpl8w6RoIKraGHUtfC5Kd4yqQFycsOigxPOMPtcPVd5EkHvFpD47QAUm2I3i6nDHNT
73knsuv8wwm5OZBdrZXvVLyZ47qvNwXR35A++b7JHLmaYNGEm574lf8ISwIyRCKPj/twH4mYrxw8
uSyH2T+lT/fEyHC1DziVKae4rCE6SxKm6E3GElgGg5jPccMKA1oXWmeKnzbCRG+69vu2f2RhPDXM
DYRZJHfdxu3IiR7UzYrZmcP6S7uhMroK1RKWwpaHpg+vGIwUEhrGsM1oSpneW1Wiu1mSHIOIIm0m
eile76ff6ozuUP+90mhQTvbrGVR5tRyUN77BQn/HUrH90WZROVFYSRr7KO0+zIiKXQAJDBjITCaS
JGQy4lnAUHt278/UQgvgKJlBgx3jm8upRy9/QEorK7/xAIJhp8Wss5unrXXZGSd4TYOe6mfvsZqO
xhQhfiMLCsEyeLN7ZOkcaDch39njjzA7JdPYE4BZMZXF+g4yKf88MalJubjUxHWKQkvYs/YIaql8
Co+VbbqekHA7JpVDVgtiUISL881rU62EYqg8aCSy/9STpZqfyPuNZUDVZRpFARXsq2g+FF/NN/UK
XjDlMft6nh2XYYTiSwiEjfw9Q2nd4XFYJ7JWlQkR1A204TvX/WHTRS7+YVt0vojN+pa6M6pHuvqs
IkpPb+xJmDjA4F1XRzEFDo1u87De/k8yVPUL5aJCNSyKburDv82JPPtncCuObopO39xiDMNN2ewu
DW1UNbdttz5fnzurGBAVBt4T60jSaGeS+pqcRe9PNN2+DHE0fWIHJgQ2fNilyVWiGXm9Oa1WTq4S
Wcc04efleT9mrdx7WYqeyjQ2icZVaAaPJzJmM9BEowInLTYoDJZ+3Hg0CSrHXgwwIgrFJxq3rhmd
NQjLQhLGvjFIz3IYbJUvSVj7h11uEJkWU9EgRz9DW51nM/Zq1dQ2HFIfgjmpFCirFQCYy0eDWKuL
moI0oGO0yX2p6Afjgo6X0lxfR5xDYX9Wxf/Dg7hViyjz9SfipiyaYw/CUTUU7OiZXxretm4x0pXQ
BSTQt7b+ViHOa6+BcaetQVyyGvPXFLE3aY7FWvN+9RbHy6WS5KwWHV6ThksiJvSORKB/eF8Zlzgv
yf0Ax84pgE5PIdWDI/ae5RPQ4DkwnsvQEKs+48eI38yZOKcNsIZ+Vac6aOoEaeGHXTuxpVxdcE/U
Ovj7hqO5X0w8IK5SXwQuft55hZXJyEj7B5mzNUz62Wze36bntyoZ3bxiT5LZqUvFulRMf585l1Xm
S8BVaRcd4dDdel0vshqQHxORDsLHUFfBYD6UngiTF+6u4RhzYUlxzvCGlHtYprNbgDKFY1vo+lj1
PPI9nULesZxHHcb59MKtZmBFcjigHCXjKQz2m+rToNhr7IiHGolf2skJHhxznvcFcIP1SyhUo7ts
OMuCCoj4CSJ6c5KdmaZH01G+v6Xhcg6lOHRgRvB8MRtJO5n+iFj2Xhvrz4WGAut/ubrhPpqketq5
/BVIUT5xpTdWHW9WJIqVhSF49yKZY+5o9zbB/afYejvP3vWJG07oy9/YEJuaEdCaPh1S5j1Rd8/c
7XWjbAPlyg4hrdDZQkqz0RlgCGf1cItlmDndEdJ7zDFG4bvvu29W3LTD2iW7bgcgRRfxXf5Mfv+f
sGnu6luXg7kUC9DtdDwtf3s5ncMlCOxCdgqY9y10ldJMotMpW5G5+Hu1lUYORumTrRugT4dUjF2r
mnLTzlmjPkqV5Fjq9hHeNWgfxChQYmUSN1zb3zDx/EGZ5uG+uV7PQXT0e2KRvkDAzzx2+J1Ik1Bd
uzWF0ynxB9K0RiNJOlhrBkN9RHcKJrkvFUzHRij6kx6dOT31RAQhLNsYI7xC7UE34UN//LGLq/OH
62vISVPC9NKFaEBR/FmBful63mY0JZ2Bvf6FhYbV8n7dd8eymYTA0HRjqlz3s7G9pA/gOhvdPovS
uOZeCfZEItnM3JA2ypGDHPbWCeaGiGHwo+b7c6cY749JujGG+kvA+PsGPghB36hvOQekAW1/vl/2
GSy/uCl2v87tE2JO2NEo8A/cl0Rykds5cZ/4JtfR+YIfW7cgrKGjCKukoWOPAyCVtc2nGr5Oxmwv
aWQAS0RyqhsRU+w/BAaA1hTVoRZK8040TipPSwFNqDOmNJ0cOvFa+DEyOlMK+hB1DsXlS817cWea
yMMMtKjGERzTukexuwUSP7LGJ1WLZQE/JN3CjZUBy/XqkBG86tbTuq+Ckq05KxIiAwsoKihtjZz3
OsUq5MGcSKKSbZ59P7A7mJiyPk+14x8eYG6xhiPLGyubJGGdGH6Z9NaLXhegIhUKrkNlNjNDxVSY
tNEfxSP1Ofcw9UIiz7xa9JLc37XSd4fEw9c+Btfd5nzDpt20TX0uIH2y1k8+7nd46543IOYTFy5p
5mSXLvabxPI3RH3JER90du+DJ0/QfUG4h/zRJsGnIk4jkKHKeL5skXEOOIjtERH2+BD51qQXfJBJ
F75INgNWn1I+2pGuyK4tR/eaYioDh/hheKoQc+iHnVWYn2gatkYMEdqEqh4t7N6rn1ek+N8biOA7
ScQ/wguUTmJq8XGxnZqacTuvMt2SFUjOvdyowKn0dEQ9Hvus43Q2T0N73pOuEYjhHtGQJ0qkaM7K
cmUucd4uZF4zSvRfKKs2g8VDw1MDFhoOJf2C79WfznckPjGsg2NvadfWXSB1DkyGytd6pcdaI7Xo
vkqIF+aece7vaUGx74ZxDcPqolOdw/F+fyhIYKH+LpjmPOUPBYvKcWmOd6UeIkOgOnB0wNrm0dNt
FYRpMryhiw2XwJiIET+jKbgJLF4bRbL7svsW49ap4NvECHr1Odu78utbLlCWNf/zxAYJUI+/uBO2
oN3SYgTQB9xAQ49vtAXThMPsy16GshdsR6It8NFEcQPDGlu29Spdz+Y8omw2PTi8tk/ZuPcdB+6a
IsF3Rl3AKCtDUAz/loK1HndY3jKfk1WfUdrzIPVeVtAfXQmsxUZ94lQ7IX8XTo/LbhY2ZmsGZKNa
OU7oOEm0NPM5w+cht1qXyQFacq3QbrS97IOw40Kadi0sHJMeB+3K+DwLvhoLZs5VQFlVh68JBrXM
Op9TWow1eud94ELAkjHYIQT9gex9gDLZ/amkE3e1lpYPMa9zB3nMtZjVKOwHK15b0gKkdZXObHbz
/N68vVujD0wy6UXtnEFLPtMAKSMdCBBz2z7or/IeKOC/PDDR7GXLXIAmEIZAFkR7/0pqJlels3du
KUNrtDHV8mpcJn+KPwXVz9cEwA0N6yovaeoI0528qytJJrjp19I3rQhlvAaIlr5gYLDm550eYI0a
bHr0i4qcrXrUIg94xnuwXa18HwSh88pwh9RQnLTvB3FO6QZUNQxcyxWD6zQwWmzbOOGQ0MJhxwps
mlVvi2QlQuaV4YOLgVhFQ8a4o7AUbAtzIjILuWKgepkEW05jJI1rtSNO8EUq8EE/7Ev0CSMATLil
KRFZW1L7bvN+kLxEIJR+Iq3RAG9BCFlbiDEBm0A7ntIPgkzPVYroR4xnn0CC1dinwdToMDb/wdmU
wmIbYsmIREpZp2Kzeyn/yD34tmQlhI2A8NgHuCw58vZQxSAkuahtYW7xy1BIdLpTXuUzS2LRdIRc
o5m1aS0FulGKHo3FlipJrW7UePsNttq/C5l1xQp6KKZTEB3xiSjVJt2SvkGOZsGiRng61+KmPccn
1jmZOO1qzDAj8IUuvbGi+AF1Z6x3kdCBdTWWAU2lcRPtSebObE60bXzxJ+272+42B8x1oC/ofGN4
2XG25cLv/9MCDX2sB2xDUIIrYPSiO8FjOSSlgGcu5Fcvh1whUvDx6OZAuS+0XbfdQfLeD6JPWbWN
iihZaZglLcI7GL5lIcBVqujZmHRujUUtdMP8BmWcyNtV5aAaJYVRB+wRStXBa6q6bZOBb2f4mjvS
9PpZlrpPwuZr3j88k23QB4GTID3XpU9BMdjYdb+YYT2Cy3jI63/jvlKm/K6CcUDg9nkWe/i4WuXB
tl2pFG0qlrBnx+p+pINqmgC+Wrqe6iI2iElJmiXk8L5uqdpta28zVrrmqbgi5e7FwIjn/PL+7q3i
JKAEaLJyrXvIMc2rANbuGt8+ZOuUS+sO6IH2qxap3q6JNBcwmA2wbXXLxSio1z3fhA4YXYOu4BNv
f1KAGRFg0T91gx4nSm50mo9RcZEuB3/E8uLWMgRQy6rBJUPXzuccDrIyPNkwNisaR75jkOceCAdm
+A7DRCPkoLQhblhSayq3Bt5T4YKEdDe+rfliDXMXZld3CzNaxfO3ZuB0h07RLiOXdPpVXHm+Ju9M
X5bcJuECEkSI5FVsNQwu1DZZCA52wYtV0xmN0H5UqFYBxwPq7DRzwevdcXXepf87Jmfv9TV3fp96
mdvydaWZPDjKagwmKhvRil++cM4LCYyXbZMfQSB1f//c2Skm5EOqUxBgGHinXRCLXkcTOHIYN2vG
t0XwJDJgaMKOC5lqpHzooaGbo/jqW8ombGlQk4Nvbffpc5tuDiQ7MRld/AYNLpteVVi7go99L05S
bYKlA6csK4JaLtey7tckBRVgEYnJie7Hsg3kCZzEmi3lT0NML2jtyTxdJtel51StBqoyadAuJxSj
erWM9nrzCtNlIQ6SdUT8B4VtdwecCMrTjp+Q40jc3wKaxwHvkwY0sFKrCZEQxFpr/BqD+jiTZIvz
K/7vRwR1j3OPZNjPWZCGFFgz0vMw6LwA1OSk2Lif4Qp/uvgDhKFKgaIuHXUfeeWSTUMkJU4i50R/
GRYuwMtUkjiGsjlto0jj/8PqPwvldpQIt1sa0MZTxqCjFruJpGGLAtCOuPdQeG/csTcou81dy2XL
xex4Gj0iXkBsMMC54mUGB96TjkrkSkkJBrrrDEalFUiyaS7iX9P3KtLYlkbbFX0Vwtp7tmW72vCF
J0BOOr7uzMmazcSwYv5u6bC7BgmTIDyj0GNkFdkG7BspchQJfDPfGEJLFNmUEmPloFRRWd1h3hiJ
OcUT067JSpQXnHdSNreQjmXxlJHix6OZFzJl7LWJ88bTpKNEnuqffdlYQmopz4ksxbaD4+I/M2D8
6lda/qD4JFx8+mUAMhHYK+RS6wjPV/SKFtdZ1vCc1WrH7rYBD+RJgODUHa6Lok1WfZUByFcEEl3M
MuUIOgyzjYW3JK13DQvGqeqHmS6Em8F4U0GEtgP5GkMKo30DbLO/3ypRq9xHmWOFWYqJcNCFkCCk
GjzO4i4Xa7tW/eQJvJrDrMxW2L5g5DpURbhIVSKe0X76D2I3OGEX4ww86U1kzL+zF3R6rXqELfgr
rxqdMuE6/fv7exxUbSJ7Gmi/11ppOX2O7CwkuQ30lMvcQ7mPM1DId5/rXFuSHpoxvCS7gvn+JYZp
c+TGh4ARvgmc7Amt1qKACvPKrPuEIXNCPlz+53gV8/VkJEGP6j9W//c9wKcsTEPqwaO+QxMsgGVB
/tr/f0M7OiT0oFKEym9mjiOQS00lesGPIw5+Bw182/vfOunI7zqF1rm0dlf1oYsaTEjLBdUPuMao
Uy3lokltSDIXGIvaenSqyrCAp6l5N28GWpQ6y3J9VGHJP7FEQvfiUgp1x+huD34JSNMR8w6WWfOv
/rjNbm+ZTpDA5HFeaB4YFKyLF1ndwS6peQ2ZNZ7N/Y6w0Rc4yUFeQBazKPjiBbmvcIMlj4OLn2qF
K9n8oh666KmBc9m9Sr0+2d25NUDf+OWe0DAjU/NffZtpn5TQw9mnzOXtZcYSzffseOu3wspmJeFP
Xc5+E8SjyitSHcr5WAC3UZcY087rotWhqu19us0vCZ5WbAWHKr+46Cj4havQWDSfVaKc0S45lF+n
Z81Vpr0rJ/5dzbTAmm/rX7GWvCWt30aX+9CxPlLyjCnPYBtuVVhyOIjKcK/Pi+91DGo/0Jl6vobm
XuZkzaDrIP4f/Lc9ufd5ec5SuENBrvawps4SnMW8oS8u9J27mqyI2MmcjQEBMWaLsDrJ2QBjJJxl
E6sKf4LCMR6DEHjctN1Au0T0u+JNU+vlBTPqEHmJ0S+XuAu3nqyIfT1Ii1XIUw1BBYsS59z+FWSy
7OK+65g6avNkcgZ+IvMCUxt/cD/FqoQD/1yHUqdKYLA0hzcoNSWnYMGr79X02TOHjiRxbtcgWP3e
Qq6nFNPZhDT7vhK32hAFK/UCrEVjOMZfm2lndh+KYViQTSOZwu2lJoePtCIHHiaD4FP/4cFpTgYB
baM+3v+Yyt2KEUtbTACM8n6hn1Gi8g2ag8v67C1jTeZf351GDK4+3KvgD49yIOw2RCqd6bhFUdNE
ykoa+YuKqv1MU4yDYH2zBndJntNNiXYC2PG2N0xlHJNYURw6VdQlMOZuw2l6DB8x998NatEwwuBu
JK4n/PuILy/+N6or9ugV33lRmQwsMBWvhQG89jIf+e4G1qU0l6gANn6/p2Rum0vhdAtKp1EIUgBD
cfaMg9rMO7qy2y78hItEiMkHsuXhx9YgufvDveuPLBJqzTHzhm9sAt1AhJwyZMZ+1HHnM6r+ZhJN
QN5QGppy0/NFi8UfhV6t2K4dhWIO9OZUxoj98vjrgsxnTJslXT3pcecwh/3taWmkREYdOsddH+wQ
gV+0cvRPmWmvXg8figXYIc8au/gKeKaIw6qGgXYzjPQa/z7L8uqZRT3zb9joazaPhX1IJfnLgUur
Dy92xQ0HWO4rYHbaqaCq/FnlE1IjFfoHozWg/toAqFue8ujIXYKTCxCkk/XuOZ0B8F+6a9J1i80f
kjgmOhfOYngtk3tC6V31TNb0suMeKDnPYbf9rghU7PMPgZjn9S6xHA+g5V+t5nmoYZ2oY+3mzfEw
/cttl6fmp9RCmsGgLIWoeF+koC64FrSnFMjVRqueyFzUPW8Wm3WBVL1TdKdZbSL3ULewqE91PUT3
TEj2ibX7lbhkpof6VJVgbzPXUECc9tvWacEgEmQq72xvTTd9OShyOt7+00tm2lRVbLH+pAIdEOqm
0Akham2qlh2oRp6WYWlyGJ3llX36CzwGCW4BN3rclcEi1YQRaBg4X5ssLfpykgmoRXG0/HjrHgaP
8CzFTf+F7DRo+s27EzDLzKuzezH8soz/bocqJsrG8r6Z9hUCpH7D7mXypj0eegevLxCKlH6dZJO3
00ur3eeENmvIgzqWoHW9MZSxWF5d2Sf1AbFKLBv8R0aMkUNXzicAbbimAL/RRbNDlc/bl2IXBfGa
C6INbM1U8Qn7SXAfHOnHtIxdMoTZRkRCPPgOcverQHwZ4Cnazsu/wPA+WamzUBbGkZwhI9yQzzo3
EUMJZ2+yeZW3d2dwcgIYauOGeSvl7UEqA9yy3lwI7UXHg7kPt28hBdg0ODUgt0EYD5C3e0UmIQpD
81VLwRIe/OB16k1Cjlqmh6ZYyjzkQPdOhfgOV2Kva8QQRJLRSmimnV58pSAH7rkNDs9gw0iZHJQ3
xF2s2Hv3TbNUOHB1bLXMZ0Ru+gMze/EhwdCsSdvzR3vA4eE2Y4b4fZMmCd1o5nTkwtZ/J5AKQ/EY
3Jz+FottwFjoXBguJPhzW89iwJRJg6rHLUedJKBiw0H0iPyOxMvqpJcShgOIs2PiVyRSd/RW+FJA
G+YH6beXAp9G1XtbL+kgq54XyRsMIJNz6y/vngPKIMM1YvrBaE1OoiapCPyyPsEg1JktykWpXM5p
40HCg2op9HDttP/KsfRtPdJJjdjqgrIJM5OjWCsYK78LQ5Vd4M526bFcBYOGAJKEwvLi2nYjSG5q
EITatfZskuKY072A8TOYzccFSMTA/Yh/dahNMByjfubub0pWgDW+EdmsLI+tQNN9mnoFNcAM9uhI
Pa5uoJgn/aFXyOvsaKliLEqWVP7csNVJNU4N3mWa2xuQRnAX2xfJCjb/jkqS5L1hoeuTgtOr51q5
i9FefDVddq1PDYlQPvallyYmbwIZGmc0o5OiLMkjdA6w27cgbPssy8xb9Rce+kTAchmaQGfuAqYe
xp5grLS3QOrv8NpIOcKTi6EziZvi5OMiCwqvVMTNg+l/OYNnZ0GDRtU94UUh+VJC7XEc15Q28n87
xChvUI3Baa5TA8VdJINaaHPqm8JBseL59L3dan4k2QF8ZhWPfYWBBC1igGGNpyWJpDdoXMZCfS91
fxslyWnb8wLaVtQo8VHra8tYNv61zlCobf2aAWkuyslUvz6eBYMv2NdO6i9jLkh28BvXiv4qPl1h
sKfVNfvqQRS0rrIQKeBoL/x6Sbzoktv5rmuOL+ZN1FduPdv+OyVv+A6KP1oLcTZb8ReFQpJYHK0b
/+qdZhVJNjU3JKhpUWMLhAgMHLlLLAepoaLT5UDY1BsTU2F4XcAHA/WaEDa0Mx4tFIO33/KisyBH
M3P3rdZMfJ8lTHEIhCzauyxdm4t9nqsuTmu4eBmi0iKiYRHdnb9yrikT2j9ORpUdW1RiNzN9xTVB
9z3eiJTbIRPtCK/iwnxGqg1fxW0mU3FFDebsFGsjY8nsw5EJ+wrznKjUg/SmlTU/dvODbEz32w5e
E23TZdp+8lwrhESWfAwBYEePXxde6kJcndAGMIe8U6w9Bm/jqftNrl8sOE/uPBpAODv/oxvF7nw8
9Ui4v341mKn6tWQAzInbpFhnI/SFrzLmB4auy5kTuYoIWUfwkq4JdtK1E1QvnIpJ/BhyhhDXDA95
3qmRixJ+plYlc76Lkcgt8um79U1tEoNf0vHDovesRnDUEqewO+rGhwvCgRkvcBubi788g+LN1cGO
e0n8b/nwJ0jzDRP36ZOY1r2fZpO3og3LWExqSPk0Za0URv2foqaOJE1Ps0b1udpN1X8qz2QMysZi
PVe/ZAgfS/cYXoHdyVypSD014JWJo+6RU6Hjp2lpJ85qdfsVaDmmIsOuTlwfdI8p5urYYM8bc4Yc
j4mFtaxs9nL8a/DzGaOEnp9ZlI4YWPUQIcZdie25Z8Yym1D7A2Mx45s3r5oWxfG01xl045eDyGP2
XZKlKe34WtaqBO2/uzzOQQpxDZ58zE4vHE3UWqn5kOd95O3B2Ko1XSZQ+jdRrRioMMsS05O6SvCA
K2dHLT9Os36J5regI+V7ij9xrdAu3ywqoOVT0MFr8SAqPdc3Sq1SCbFI7eBtGmdMheMV0GFnxoRo
6dv2+o6iEJHvGrIriI9M5TfB3DUps3/3RHSSQRvigf3dWhNhEKdstX+XOMZ96Pyol8XWcpuEVbgr
pe44p/QcHIW8xKHwOAG6bWF70P8YSDGqD/LHoxE1pvdjZI3nE7P/DdQfkjt7IyJWYZlsAmpt0xey
nnAzLM3d/W3hzheOHXW3T6sv0FhGQyxaMBHWxkM+M/UQ9eTMUf72WgyP0MHj+r97vRgQ5Q6RcxRi
XU4R9UjcYpz5fHlGtNtbMcjlOYo/ANPpSg8H2Qgs9IQCLkFTLiqB23kRyub8LY1TM/pOenxoW8iF
YLof9C6fx5l84DlHFHlvIkYojRc3eU8d5FI3JWw4ahiqPdhZA/l4A4R5pBgxMtWNTDjWhm0NGJ2l
eexobMwv1kuQhVlII+yBJnxhfu9UxzE2lO7BIhcGhGHb+RaNbfo9GvrErhmLC11Cc4/I0sIUGsMT
+Y7MaXMGR+lot4M3jF4LiLO0CH42/mrB4Krcod1lpdjz7mwl4PKdPyre7O3dmm3By0YTh5dchLXU
ypVI4a+D5+02fMdTELh4PfFd8N34fELAopbbfsKhpZK4xd/w1DI9iiAUdWD27CZamuXth1yy5JLD
CaH7N9K1LoxgPlHPzP0ze8dT0YPXamkV9ErEaWMqa+OB59HoSdTSXRjMKig3gmfwJUTeOe8Y7oSu
7QdtWlCV2TEXMpzQolc18Z8PXgyaqCOORMHh4rcT+emGRL3lxzd0XMwFOfBbaj2893q7Ydm3xZdi
kuZSV2P02iLsW8YqjXFSRE/WJ1rADIiR0i9xFfCYeFCc2645XquxufYWBy6ZE6H7uYZ7dunHTWBd
nLAeAFMouv+AXMibpagTiMr33tkSCi7G3sFojrBX/Lchl+Et0NmEFgExhlP5cwJUnIY7Ha+IrRvg
KF6cHDy85Wf+S3ddFrLurj4Cj6LIvom9TOYic9v/XEVT7qGLrvMQQT45hOabN9WZZBctnFyJWSSc
zMUEJ6bNqL6QIppZ0t4IIkNqm+Gm4K0yuz3iYHxVwZ0j587MmETfwP1WFBe4NEWG5VbkiGrnrNrQ
/VXuHn9bjNMZCZQxGBQkl9OPR2KmawT3/RXjyg1uExvIJn4ZcEQXBS1FDXL05jpFZODzTPQgnmt5
zWH6CcUE7V4olbJoBQmaEKBVoc3BvdiuY2t00O9w7gGlfDapw0fN0wvYPKHa+Pak6qpAMgelUfRF
rzFwJDW8wGyO+AEkNmqD4+h6DTRpdZCJIAd4GH/1hdjMKvkPvyiN2UMOhjyr5BvNfQObSG8715/e
cbOQtbxPu2Gj6Kw8oTGmufTosJ5YOjK4WWhurIidx+mhVB26aM/0fIs2b3bTdboL4wcoRcqTlt/u
HT2MMOY9++z6uma7weEhhstz+Ac4+1vhEQ+5KZoK+WxlXdUq446DdUvu9NUp0YQ2iHlrnvzxrX1E
kP/4pi1OJT8D+B4Y/QyEjiP3evS2I3ar9RPdq30HRBsk6qIMdr0w7TqcZ9MAs45qPnS0WEKQ4+Wf
tckW0StU58yG3rJdQKjNbUVMK3FaAs6OhkcH0hYb42b1X98839d2lq5WymVy+qnJ7s9UwvVET0tH
cHhZC/bKe2xyGss/0FOYkKDdYt8PSS8eprOnz5dGgOMpttgByc13TLLvGz8JU71tdhqu5sVffn4R
x+1QNxvOAem0UwoznMChiB3SP1TLIhQBT0Wj6Ib6rYPSTe12R4vSHuaG0CylV/nUg7J+W6+h5Kyr
GsfSGCKYH+PX/p3HI2AUQgxZStdXCkIy46ZPvLjtTWwo3PUcZlj/BTXgY63Ekl6qQiFq0qefRy0j
waPlEHyseauNPzigDHRtIVk61Sz9ALDWJjQ5UDYcck+gNWdtK661OYrRxecF0YTP1VG2IZGg8Sai
62lgUl1JK0GDzeCnsriO14kqir2ocbN4bZwc1GcK7k9pbpmZoQCfuppAhMpRa0fpKAPAS1/I1Ddb
48mh+9YaLqUj3rwTkY7O5QDUomHjL2/MygdBsLVNtXSWSseM2Nz73gK/yRFjS4epQ1qHT2GNszBI
wvCAzRevpGPpQRx2HED0MOrpEDy2Z8vyKrRSuAbNu+VoGmjMbQwLBi0xQj/h6H+Gpfej5U4gFC8Y
a25smxU5gyLCph++vPzLpG8/0WcTlmbBNQXJkYS3nsvpXIaWov+II16ZXWcgm+EbJi6s30vLybir
8ndDbYUtBLaNAQ4wBzd0as9derH8j/RURETyN5q3p3euI/KZRtPJNr+tC1dfJ5dTPCKoDnCs8F0a
0xBHto/MO2SNXwffhHdIaOszSrXY8J8Hb8H1cx57wo+CPvCXVSy4GR5bDyAGF0fTT0Jl5uBtj8BV
CLKabMABBgjr56lNIAkbdLu86RGPY7fwvQO9T6RsiBQ1y09xBXuehjP61HIzYMK4Qt+xxVIrqAtF
wFNKLzodu0qUF/95TTp1oT/jhTob7grZvxbfUGYGWaB4sc6fPU0Sq8LYJ9tAblTS+okOdIfzf+OI
BIZGB0j1ER5QHYTGQ5Qje1SLQcalKKtpKYTLfBJ8qgu9mKvkAsrRpTOMQ9+G60Xl4Yk67dCVWGMD
dhDXs6Dom/+yr5KzKeGazykBz8l43grClweEAzceuBi+C9T1q+UPj4ugJ+jsmACIe3f2OYUwz68F
IG/epg5KkMb0j7qgknQw64VGIkc2yQuiEGWQhc9yv6VMAe0zV8TlXtjnksmhRsjpzKZiJbHPstKV
NC83HwMoJ9ihppPuSH+3RYcUd8VALn1FLmFxOnTHISVJ+0Gb+TxsA45GYKyUN7pkGOjtlBUSyoLB
n/mKx7mkMl2vQ7oioY5rF2miZYHL/PsBJSaBETkcZXIWdfiZXYWBHVtAOd/LWjNCrPOTw+nCbcBk
nG1weYCe47G9+Ei1Zm4cEfcADDjqheTrDLfYZtXxU8tD69yDUGlSKQVTmvpfRgnyR4fTs5H5FCXu
ivszk8GHQcWjKe5jd/O7ECmgisf785UwuTe9qepTsiqLwMbjYlquRLU5nWdCmFDvQMhCB92avj2W
xXQQCH2LX8s8DFG1YTPImov634+BkYYa5um8RTLBi5T1wrDMhYibppz7ih0teiKCq9P2IMvLEI0I
OhKMAWHWKyP5i0SOqkK4HD/Ss+y/wdj8+/ikMStjaXroGO13TmyemThf0h+944I/eETpKS4cFVVf
JHiMwuP+o8xxhJaKmGP68E5qgUvLIILE2RMqrQBj8lLgD/3NyO4s6uZMnjyRCDB5Yf+k1aUFWVOJ
6vv2YmluaJ5nxpbCZtvNMSt2Yse40HBMeci1xHPelBQMki+dnjUuNu9ZKOH6XN6xwxLgsjcOrlSa
ffQ12aAiQ1LmN9JFNhBMOzDvvtM/mM7AWt4/xm/teoESVLAF2taBxkPDnKVabSbYFvRJUOfgV2qK
y1zOsCJFKF3O/037EWpM26eWjSrAer1PlazqdfKCpenOn2aSZlokkOeYLlg2W1iNT5eIgj+m+NSW
w8cCvy5b5YWs+olpQ14ezZcpgmQzjzc40vwscvhtuKhEqcxV/a/0Lsl0Ym50iyAVbQ7eosUS+o4o
8vUFM7ZVRrfjdGDJMFebq3KxG6ej0Dc/UPABprLMDVXMFMDKX0iJ/zm+kojozQvUIErPQe8tAVNl
Ue5i0g6ffICDsWqXtNFxBDR7EJoPTKuXbh5IFqIwIjJG9Q39a1TZJP+r8oVHg8Y+iq46w2O1rp0C
EiePT8SNkngWkThxoq2tGNofwZI5wk7kf8n4U9O2teNfJsc9sL1GCvm3TdPQdPdb/AmfVarpnHze
Kt/LWMESW0ioXtl4YIspD6AlnOj38DCcG6AW4kPSSlzclfsw9YvN4Ivi/px87b9P3U+TQZy078OZ
2d5DMIsVBivCCSkJliJotsKfqs4UWEhDb1cBDUitLHRJ63DMu5KWQ1qskyKDdJfsySQQ9VmUEM5K
Vdlbx5URU4a2eIgAXyGg1xRY0PHNBPYyt4eCnJkXE8Wta1E/Rfoj8L5G4PL+I/97wFueVAw4RSJZ
yvXH8s9JTepRPA24iPC+HnKtqwkLYDu5Vg8fsgWY+N5rU1BMVbDbu/i5slR3RA6S2M7HScq0baEE
mzBTs9RU0hBz1919yYDc3meh1msSRZzd1JYtz8U1nF4nNZ6sPcQICvBJvxMAFfVh1Wf/uR+IsOoo
iN5utTWnnG//RspRouUnI+ZINoRS8w5ECY+r3IABpGBCRlGx4POd1mLMAbKT8d/QcfLPEHzZi2gj
DCV2Kxvh4eYbgbQ4r54a/mRpJkumaJKbpVFMiZQ7XcMUWFuznBAsdTfSWWjXes5m5mypWxp9IKUq
lX/NgSWhXdfJndAaU0x1m8N5o6Wjdev6/1dNnEJgVKnt9p2M9b97VpYPUFVlPmMTXC5W7bx+dQKY
AADkJCH5cI4shwYZ38YjfZipX4NlyQ6Jm7wfK1KXuHE28nPp3HOP8Rdp01XqxvKmKppIdIAaeDzh
sHBzHFakb4+3BupYzLkIdyQVa+fI1YZp6wKrzqWhG+8Fu2TdqLObDuv4HR06DMZqIFl2whsD6xQ7
itvc9+tyQ/de+Lg4x8HTBvSa9cPoIdlTRkZWSZAtE2FTe9JX0eXHewRYKNCMgRg4r9KXy0tZt+5W
tSp/s3h01Ll2AcMUucupB/DdmKRbHcyXEooj9+JTUyydkwPsDS42IIPgZdZRRHFSyC53BkTwlv8N
sOioK1YGjoKdlG8qMAgG12myTHrXVqnBvmkHbuO3rlABvGGMu0BsLXLJZZjn9ZMLobtXtEjjUtyi
uT3o+tUZNrjEoI8azrYfA0JJK1u0buSrsoLfbmMSs4dbruk/lqzYdMITb8pz/z2p071kIVeYTGMg
4lJmMzuZlgk0b5eoC3xJzNb3s6qrXkmql0DIWGLCFxxbnjSUzWimcYU+A+eSDioBaUYYb4wVl6Ak
GrYt4Tq0hQnNggVdSPvgeAChzje98d9MmWWQMaCRcN9pCIc0hmKR8AR7v9m2qlqUkRraEoVxZAhT
KHKczhT020RU6OMPwQS3HVpYS/ukihk5deDKpbIIvsy0vp9X2X21dDQvkm/CfFS/czQiWnvYrWXE
Qrg3HvgHdoUz3i4aVSKMmw/7lACQmDH19ojjJwOJzBceA2wvGwnkJDx0hjc4ZTdfey8F0zYcExkR
qk7/G7T+efFUS4L0jUogJ79BL7HiIuk3eCad6ske3aSIzRTeEG7hqZhfMBc+zHr3f669mg6So537
acNl4T2fOnVnJxjbhuxQawhOr/Bq8iVYhkxsEdRucwamQdzXZ5RkeXLiHrGnycHkhrS527ruPuuV
rjqd3ci6iPI4Qeyv1unDk2YAOXWnRL1CBfnYy6+gLL4tK+yRGHp0MeRhXZr0F/7GvXfp9tlQYNLb
NQf30QB3sOGBiqGamsFsECJl0v3l2xWYlpW9UPvf7tq0oFPcYVwcEicOc4/J9hGLgxIeKYG/8TCM
PHlOfQZMf7iEQNTLS/M9VpCrAHOBFBlciU5GPEIh+XPpWd9YEIB49I8IXbPYBunC0YitKcpkxtRs
fAwz/TBBLa3NK1jcPeJgw8cVMbdbgPH3H6LaqPDkrJEXvyp1DFUViyeZBUeo7N8qe1jBWngLaidh
u+Erza54KhnFykMhQXtECC6eqr7CAhNfWXwT9VzcmaXJEBfvrEksOCbGMr+6ctSBRlgDOe79F1Qy
t8J3qxhjM45ogRrLUzRjnDuipE6WOOZqsgsvJVqUVq5ApSX7dC+lIgVc+ubJ76GNZP1ReQfTGbNa
2f3XfI1IFXPOh6o/3w/6Elej/eM99vUhPQNE2cU+cephpPRrcgOg76o6PAkurYYaec84mQ3oUSrw
I7Sg7EMdWt1Ef7NCwsEzbV4ZeHq3t/0WWNHIE5e9wqGYXSO2i9gTe11MgCGQGlmYxaJz+GynzpzR
kNgB99IXTTiLCklLkUpG5MW3xOMg+w+6eXdL/lGlLwIoMx5MhdBtFeBokDx9S9POQnbOd2cnySnM
+gXEK5H/rFF4XA9FV852Q0HgQnKiuCT+1pgPPuCzjGCrFarvzlrp9eL4geYoVwHUTjorVzM6K1Cj
QLbrXJ9bhajYqn+AiTjqNPz3Gv0UYGa4Sm88PGp+HKyuWp1Thz7/+7f/ZRtJuqSSlKglmf7FAYHm
nrUvGPbbVrLrkyv2THcXaZZ6z5K3JeEI6UJISt2yqooMdw1E4aCHDsOWvY1DLEvnbMzIZqqEtNCt
OUKJZCGSa7i2ZGl2FV5PeOULuVwjUwnk/PSbEriKONeO35PMOQgIAdyuq2KaKNLd+ga5ULu6ZNHk
rhX2Gl3UyyeM1+lp0svFjJhT9Sjyly1ql6XxpZo5TV9WazlcEE8n43psE8cgg07qOa8jRw3gYedL
Ejs6jR/roiDXxir9HHl0WREsVTNvksAlyXmn6uqnCNJCAOjStopE4DNHGHsG8EmICqMvbLv1pNu8
4UwxXRwX7JmSv8I+YQblkpq4HvkSZurSBOVVSkNIUCvIR8lUaO82O2Vsy+eSXjiLaUbtrTi8LZqi
IKeNndhUGYDRBGt2z7L8vYcgRRx+fN+Du0vdKQ/1q0LKwSSjwvczUHQSFcR+i7Q6JsLZQ2EHk1c+
lGjUwBzdr0VkZfnsHxVDMmAO8ZN+D4gSfzPjd0UFascW2ezjjHKatMuu6e5UrrTHbN/8st6W5ilK
g4Tu1QICKbr/eWHL+YXf2y9TtiwKNhcAbfjgJsasOuTbSI8rS40MWcCrjD7/bCAurvZTLITsUb5B
uMXs8rRdih5KYsf/arGra0Es7Tvaas7/K/gVj+ZNGYler1y3QtBFXfnWIcOXj6XHb1CYLeWxpRN0
WmDo02wjPUknOaKML3Hjt9Ay8bi68Jes6X/nXoNjT10xq++NNV6FG2560OrCFxvXog1pErkKuhFT
pz5Nzbfv39I6Zp2NjsU9anRpmyfPKRQR31aDlER8Vi4YAuU2/N+esp2C4/xsxERvHUKJz1AQ66AX
r4dFyN8iVbeakS+riqXyqI1seDV3/FZxmLlmR1cNT45gnBK2o8Giz08vqbjn2H/HhxIZsKfFkvml
wPBZcoVXhK47YFsgmGGAnJB/v6lRGZLeb8omh7Fi35c3kDhi+RpF+yoahLGZD4oZJngAOyZREwI1
wtD6NkSRPZPMlB4FgZ1SZ+vdoWVNcMh0CxpDwg7hUvUm3Svr+2KJvoJrdgjpQsCtQKWM+V8LkMWP
iEUVTgGHnpSklX81bdCIhn4DGaRHSrmSknzciMzzsJSy05x2utGL0NwAzLRTp6fR1SZm06Z1SIsr
Nhtqc6xvMrANRbFwsDvkIQjxqelA1AXYlJZyyWuT7gNkE+5a+dE1QeNG556CoX96KlE85mEm1d9o
8gILB9/VaBX3+OnQQWP52hDd5UAPhnjB+PjiwASoSR2QNVMR9XekLCa/H5G+svUOTXs5ZekTULTV
C5akMcQ1K+3EhGliKSIcGcC+C5tGSilC5W1SES2dWDa0TQRsF61AlZrTJ2Tqq1+l+qhH0tR6Umh3
KcTG1toitv0u4ieXZ0+eGbtLsA/xVwniX604z1G05QR+YkbL6YwJtwXEyeOC+l2jKDrxuE5wjaM3
8o8ZhwL57X43fkwruyfAZAOi8aNHpKo7wbjKn09/cGte1R3tAxmGZMTPHn2CfCEOpKDS5UHkJvqb
6C0tjTTvZQYWNiLNxT2YTBRlhSc6wq4BFr8p8Kd4n+KyLvByQzMsGCn8xE/tIr9zGxkkTnlTldPY
O4ncbDGnyHc5UnE6meJYKFn4BWZituGUq0q6gbRZyMsH06hHkVZUxdUyx6dmNsFIPDzrXZFEoDLu
FtGqo4+RqTflZNhNJd+S/Nh6FAd8ysz6pZ/qMRugWOU1EH07KV7e7oc3los05z2IPSA930xHuzPt
zZr4RSI0ImJzDLc0oGrmIwhA8adg16Dx/ybC9cJ7XLqCe3/euvVPwydReSnh7bcN0JxSZ2PycVCj
Z20yQAOl/X8+V7c8FWe4uF2sb6HVvoj1UIhP9YX6j3sfkb/x5gg24735rkQ7FPSFUzrLJLr14tdz
If3inVzqX7vBk2S5QDLwPytSeKamMxmj7IwAmfNcW0SmZPxxECM9JWGDZa+12EK8LaF2q4PBK17s
mus+SRMPGcyCXExXMaTG3KLS2q4i6Vl7ffk7uTaQ5CN7L0wtYZwsvcvd41J/whuBUg3eg/ipDzLB
x1gIHhInr+1nvQ+S98mix0KUCb01lXdBat0TusU6RWChkzeSY5WnPmk3xgN/VuV+c1hYOSABnHak
dbJ0VPkaOVLiYz2AD4U+99nabgDAljGQ9dQr4/72UzEX5I2oB6aVNRh7QkbbEunvzW8pVBvVSiKW
lCKPl2VmODsJFAaw65stWUWIrUkLEcihx0u3CgBurJGoBTmnVMNQWaeOzSSOvWDb/D0HPBIlHrjR
ITzgtYiMP1Gi07g5x7wzKm8JGPf5rlpODdzv8EzMEbDiIeP0nGrLTtAR0efLHQWb+xWGxysHqSfQ
zyvbhZ5A/ey7mz6ElNHytVzFimGWITQRKbl9K5V3mjAajzmZbADjmFAr1YmVn6gV5B9g6UxOT0oO
JWblauetW2VhB+XXYYwb3zSNKoq+DXv4RUUjElF1VP5WsP/9CoOfItKehAluYV1/a5jQujz92g1N
TL5XiXGBFM/gj3VApYoPGJwZzx2xGdWz+rDSft6osQ1XwS0WQKpnaB3DGPY4grGdg3rABWW5HPAR
0/JdYa3z5DaDKf7JxWQlf723lyOjPp92IiXHGBbLuf0ZwEOjthncYfxstU0iytXtc4LlTdIiJNvN
yrIoUOZk58UetnKbJs1Cnj3N8UmfHTOkBL+hkqbd4bYMgmzEpA9dl0HaKCZZUjeY6MaM7RWDZW9C
tgQxM0Put93lxKK/uPMKSBoIZAl6R4vNgoYwYGDMT7Mlp2NvDukp5fGKQAtyAwdFicS4w7FP784u
LSBG9mwV9GvoFCgclfd0CewatJEVc2BUAVCEctYM5CBVu5sdLQl+Ubw11d4fjyh9AAnybBcCVME6
FyE+HkgqP542I7uUQ2CkOum09PAZnCnZlp8Lg779DqsW9rScpbRz8RndkOQX4dmwzUoBiYpdboDA
Y0myuezfJBwHYbsUUBtqieATatZyivl3nE0r4oct9PPwRfx1aj7+5FAyihKKPgwxpplQvN4V2JUs
zrk2rS5/aZFrzQjGd7FJzJQq7Fx5rcMMNedL1cFy5Asgz9yc+vLUYwosna8TNDo+dzgPINWjST4+
dAPQ04HzKq9wKvAbMO9jtH3ay6AJbcV7FXLOh9NMnIegoQJjgcNUhKcT7rDmV4APRA9SGr/qOZvZ
l1UMxPZ6EnojVwpxrmkIrdyR23f1El94vCtw/oJ+DnLo+JH/PtrbbPO8dx/FhNLTx/lDXjG+Mdqy
fWUOJavJAzvlySjlfTvo1iddtMJHzOjmpnmLNmu0a0o2amRHqQjgfRULPHJR8+L/56KPMGfiLxgV
EYzlTTxVIDsfqXzOldEQHiq5P7/nIAGZDPV4nNM71/gh0Bkm8rQhmvUvY8UOQrqukYlLaMa84NLN
ILsjL28cS5voFaJB2mbvb9Kj8eqf4rbugdiblDyF1ZvZH4beSt7dUg86TDoA/10FlI2wrE1BIlpB
BzW3bazbTvNrtwrVyNsuAGikHiYb/8hj3QENHzG0BNOgfks6QLpBMewt98AfTYitl94OnQ8tbAc8
JhR+1GjdxU8HAE0fKzfdMG3I4bsUSdqFNYveOs1Wp83Nx3dg+E/qbbkbbFpK5C3lrddvEcZSXiF/
1Yg9FvvbCROmVZiVWHf5R8ntPPpd/seTo6MCl697Y3Al+rxp68KJVmSk4e3mkmIR+nviryOXdMOn
JIIKYHoatxqZJE9sR3N6ceBPlqICJLYZ4pTryiUrboN7ychqYtrafElvBj7iiIJRBLkpWLULIHQi
p6mWIB9GArXGf36tBnP/lU75BhceHQTfqD2aOd6rVYPYEc+iej2vLF/6xIZHe6aGiC4MCrQ6E9JE
WeW/TviQ769FlcBljvOiNt3MJMDyvCGKSmjG2kvnv/jEK+QzvmGrmATIxZvmQPQ6zi2AgcrDjUcu
LPUIbT07yIEL4W/S+lEnRpKqOJZnqaTyR9OSDjdARXJrSOSIcQhuUOVJ2bBPmYrxnqD6ggUo0i6V
itVfaF0JaVCaxsVjZfJpcl9evBN6LWZ3WUeJu3ZmG0GaPZ+ldvoqzDGwL+sbDDMJsl3IX10z4yVv
D1lFZmwP8K1YkgLBOqIy0P28pavFbGVdGhYvhI2xcj4Ssqpp/41XSIme4cQUmiWXdQYDubrJ8uWN
9Lwfhb0OhCOEaE9Eb2XFyTfe7cLNM+1rwvm185Y6RGpWjoZkaVDjsGE/Ic3qD6xxq2Ta7An6gTRN
erc55Hi9sxny2FOhLTiWb/k4po8QE5JYalFbzAh/q1245U8Itc9xS5r89lnkML/I1G4ed+XOBhzp
41mNg2e2mViF3HLeEtCGsQBWdzMLgA/LkLKdixFwAdnf82zRq/wejpEPt98JjmPBK/aA7Mr41wWl
9zb9l2P8uU3zFrpaKxMvcoayyLUYHn7kpKmFCQFE+V0Vvix80juGKXGZRO2WwKwRvi66Mf4sOXCY
sEeWcEpjMxD+V+r7gzcDbT/NF/yMiiWee4DsPpmkLuQ6BFh2HKfLKPbP8N995Fy0E7oUT6eHqN15
n/F53YABuY3jGvTKL7S8jMU9NhvLb+pT3kDxNZ0by4OW7bSPRuRurAP+xnlWf36tLz1wmhDGkyYd
xdTf3ebhlXa6KmfPlyNFTKcnKAHg9zI0XNpN5cGK8J+Sqn3Ya4JE2J/kwTOIAvyIBxzqVJgt00qK
EY5rO/HnDJILJFH8Yxv9s7FXI/jiccM6ACUFbL6XC15oL/eH0fAcb3yTPK1tSTIJZGNFCLMxqi0+
bfi4TTXDJo0md1Ro1DTuegHCvmPbWNiYs2pxTf6RqhQyfOHDfxRUKpByD2VM9G/z7YQ0h5bPArG/
9EaakEBY3OlG1GmHxz260kNvNK35IHRNwInWkuXEvTwnUKNAWt53jTICJgFdUmgqr7byIQOcfzqr
2UJaFKS4G3aWELQVrFUXBELa7HmAemmS47evSZ5Ewz85pg6wgh8Jp1noWl8GaFa8prs0ZbMIgxTb
WliMKzIaayBbtsbVHdpP+u4iWK7C8GOC4+dNwhsQeF1WO5PX0BodZSRHR89sATpxlVwu9k9hARSU
gLoa/aq60XNQNwQuLuhDDFTHArehEr5VdvprJ10S+awIHM/fy4tviJ2nRW3PAn53NM/WbwtRC3oK
w+X9hlv9SGCqeUkTZvWiTGxFUrvnE8PnhXd4UFadkZPQYzFiR+ccyh0dbY66R1MSOpzqoaWgoBF+
15y1nKDOMxwb8qGZuocStVFTn4r7RMoKP5lUfdpfrs7uK5AA7K48+R0QFkoESfrpCifBrmsj+mnN
KeJ6D35X2zwxHaianigm89PA84GUeEeaJE6MJKiU83DPycimcO7HYnRHkRQK/V/2a5j881xJH7HF
s1B3qo0yNTgmo9sk1dShE160zV2vS77ca1wgKa1+tSCXsjBJXwk0NBDH24jWhRt1K3RafDlAn1M2
PDgncWOksCtGX/BGeD5FTZlPTRVyswNCyCNZWX7JxKTC+e6LA4F/7/eGJ9Ev3UPmQTKTnZSmywNO
DJCHw6DT92OCl8e1BbEuw2naOI+LGag1pVBkC9XHLCxCEkggFtUyylPe0cuNYyRPlFnT+RjYlvfO
ohuD1ASEmwHmGhu7d4Z6vP2/FK9CgJRiNVQftTIYUGKd28jF8OhS5tAerwg/XcJKLZFHJVJ1oGCI
7+DUq2xpjBpLKSTzKSWvEn6gIPT/Vkqf8W0BtqkNVDgrDZt9D93CrO2bcKPSrCxUENp76Wrv9ibm
Nkj1wctiLJXLdIFgqOTEKjVC6VCN5rmOJ5Ay2orPqV5nH2oaTeAK0QDbaqMahdq1fEuyaURNVWWI
1O+797SRmOIcWhuWDM73XAqBeTHGi4/poyTnd7Yt06Pmmyhm6zsQ84nIK9YHh3L55NfG4D59o8J3
7Z8NSTYtfJ4i45GqoaaRA3VrFv08ET9Y9ATp5yUo/YoVfSnW1VW49xqZZx6QUtrn2mwOFtGlH18c
x/ipXbKM56/wqftoBPcTxGEVkZnxkCFFsC4DUAoUF9CcPKIda/d/C2qVedJGMQQHT7QAqyWwaCr/
xkFARBoW9xINmG4LD5/LvOD38c8XMpu3eNMwNMx8ybuGmtApaiKi684WbS9Md628rGfOq5lpxXqX
WqQoV+fRXztuKAy7d+fNEL3asZXxkJvj5v40j+Y5JSXUoYmhdQj0Re0qYp8teH8htG5OkkUs4eTF
QY43ZeaNySR6RshqWixZCPOcTlRI0AU8rNuUr0cVTVI+LNdsd64PR5RtHcwiakebOxGnwhqLI9eU
ZTlK3JqskjaGxAYhuHTPum32dkcwB2wuzlkHvKppYrmvy9Z3fk8oDQo/wtO4XWKQjjM/KNmdJMPX
h3rIZRFFvgdVnk8ZWi1d/iY3r1jU4k8wTNRihETMFHDK3XaOAo74diiXNIvGoKx+mMjmshE/RD3S
rhN85Bs5HXsBT71//d4XOp+MdxDCJ96yELBWcadoEwsSs+9iPECymxXXrI0y0iNj3qIDixHL//4Q
S1yFM9JoffL9mlGnC2ITgR+8dm5wAZKZhWDVS49vgvStqAQ/wVxKqiEd4CoQh9tfbkCikSrMlTEU
NYHxKabaPkGfnHYEumfnsBJQjr/Yn8kWtw8VqSG2zB7lp1fiC0QZ/SG7vebnqu5V9Wx6tjj08xqu
aBPshKRqjhxdPo8uMwC2ZfUXu8bTKMtH3bn9Exy3nhSmAtK6Nxd2Vis0AT2bDPqMmwvr0pM/j9+e
FyfFZajdsfXmWCjhKlyEIBpLRBEB0rENZplRejRE77WdRc3KVsvEJHo2Ef2+CMJaQMsZPOkWF9gi
BsYIEfGILcCS8SUwAYyPejJAzDoOJ0ab1Bdq4s0G/JJtbZUvHXpWYPvme34hExV7VM6bOPwuRP09
On9oGr093H8ayk2sNAVp2lTrAby+3f1eb5j7MjVt9T0KmoVLqjvUh2bsAzk1unD3GiV85kQZmi9H
gwn75MRpSdUc7uzesLO89Nm9UDlCPVNxre1LG3zVfo2kQnfHA01F0H3V8XHfRtplCO5GPx1w4upQ
8w6y7kWuLrkIb8Nd7kSqzCKJ+vtjRDBRMAZjqgThjtK7/QzD9x8HsJ4ZK0xyV8oTzQF4Ji8TMkz8
ABJc2c5h6d3A7noccAoVIRx49Zb3xCdP2MEvXFAp28kfk2iaxT54dpz7BSEncXJQUZlpeoK1sZh9
NPxvwPE0b7ktIVzpwoI/Asxk2OlzaYfe2dvKOLtZL104l3xZ0ZMnwIpPhoTXZ2Kynu40Fa2TpPpk
V4PhjJ6kFfBGtsnWhUjwgWghCCGUsuXbvg7kI8wzy9KdVtfR2kAOsQ2A7rV9AbmmhtA/iFdBpbeq
PmZpZlflkXAIYmLWVyFeV34m5fWvQ1yarxlmDa8rGOcvFs4MJmOoZrrM02nrr+v2xOOJ5qsJqa5N
oWv1l0QUtJzr6Fs6N8clg26F+my6u/vsa0qWBGTjAtyBLfUanVbtjtYRfy8tVttwMRWRciiGho4X
M8gefZLnLbdlSJaor4RVOUfX7O0VoKLsk+gSybPCP0J/qSwCbZut2vB2AzujxYQ6emlCvXGxlzcZ
V98IkgAbEpswLoN5mN3oSDikRHRaP1lUY6ZHQ65NccNKcWHYiOA2/q/gTf8O9YtbE0tjygjctyy5
xFS2mateu5n1xmLde84K4GECT69XOqbFVsjzl/zKobKE+f5WQnWHBA9Er9rHqI5T/j4fs5OMANYf
rR5BU/Vet+AV3l8fVRp0L2q5aml8csn420ngkRLDjyD482oK/ojHSDKyZJLCgvoU6N9qRQD/Ri9f
zIGf5xv1IchTk2DB8Vz8utw6gUrQkg65LncNTepmlYfOvmAYmBUwlgcmEA1AQC0GblYBatBlBzwn
oMiUH+xDSZpguXWccNvROJJfaS9OPcXH4IGJ6C5Upwy+2lVeApjfcxCpLAWzND95tIBo8H11rTqF
N0qbH+DGlheFX/Md3ZCJOn175OY/gjYiKxCG6yGQLBsgjggQ85NP/kY84m8YxKv5sYmxGDqUL4Es
JV+ThA1iqB6FszTV04KvzmrwiEOGJUWL+GNl+cYDwsmofTkpoaz0IjPH9XQ7guVjEWxBRBPFz3ef
Mi+sj+LYuJJMMRH0L1/tgjXP7I/2Bx85+RU/bOMmLnGTwKxGnaWZSeqCL9MW6dHYu/7/yMYB7Jgc
OCSZ1DRj+e36T5sQ2A/TMmU+xS1bRjf/jiYf/EAOOLH1pzPr9UI+JyqIIk04SG8E7XM/D5/QBM0j
RtVecePyX/IY4P3+63vYl9cvH4N01P0DYeJALF6oE3AezlSev4PHZayA6Ipa6W/Vbwjs4uEZqrYB
8XE5Tzfurl8ZrY2GcqpLX2J16R5HxWOxL17HqjLNt03itzqLGX5ImN0rLJ4lGPbEk3fR8vL7HrN+
LkbFMzy+MFsLdBBmh+Qk/Q7oeBCKyP7RFgCz3PWUaj2ON+de0kz+uA7VdS27yB5CbkCGSf6lkuvG
xT7E9fLy15prTJ/oTdSqxZF7/zIrz1gxB7fGFEkQ+0dW6mVSG7n8CAKzRD0SBuJ2+OhlxP/c+Fzy
USgbj7iv9dJjFMMrL01h2ZwgCdWVtDOciI3V7mWihzFAPZWjfXrcRx9mCnsYGGwRLVAlbdKNK5eB
00E+jPKfOjTpG3JqUJe9R4M6uDuHDkVztHQXjR0VaDSXVUQD/Ds8ZnbJuHDu4ZejZhBfckvLkCIU
qpBkqMDjI3MmxfiQCODJobbXYvo0trJmRev8+RszncYMQBAe3GUJPe03mH18Er5/CIE/PVng7n+G
iXyTn9Tr5NEVFpXfoe8fNWWSGWm4MzR3pTBLKBCdpGtAls7efa9EhEAPi0FuSEGtqqdorhZ6HqMa
TjFK7dlNN2VpfKC7Viu+C29H9VIHQg4recaVH8VOfvUUMp/IBmeB+8JlE0PvfHfBDqFvELpucJ4F
DMvX6J1tFT+3YvD8ZjzHuk10+7PHOgWB696kwje6DHJBGsYEOhAHMa9+B+waZ/1j7G+o55HyORM/
rBeEmzGilkutkHIsCZWf1A4saoJl3RN/ndpCrLoHkXv5YkKVrskS2WP3Jz0hxh6XKkNBI+xDui3G
kkVPiHEw9OxKXFwkvZzlh2ehPq04nGfXlhKFMYWzP3KiJjGmlz/6ErOXTA0gkPxZigdjOr0JUk/8
lLqMmG/26zvRcQrbJnOO0ge0QCeeDiNICuCM/eFlMYcAn4tqvZ+cj5t5WsOOanP9JlOgYRhWZFkr
Az1+OvCHTSupJsmO1mnJ3CHduqmgOfSCxcZ2QQiHoGb4Hs45KGsiu/eD/JBav3JF+WANVp2xGsvl
CUzfnKxcY2WA9CwfU0Fvtesg/66i6ZMTILzYo+nbr4/AOrGpmxUlON2r5TfKtMCyawDqh/7JHqPa
C1ka+2H0B/TS96xHfGrx7Wmcjy2yYGCi/6AjoETzn4t/jw7ia1KZi025lnIu82j9/tH/88meA8KZ
Qb/fW3bbnBYMOTllmq/TARYapouohD5K0X9MOjC8BpXCcym1CpzSHD1p9X91dUtJRgcrfsTv5bod
wuOK5jF/JcLRY2w8HazOOeUjBnrrUEqjMhi8kfPvFpSW5Mv96Il0ZuqzWHf+bvO19KYHI5DnRaYf
xfgTEHpaxpQDdFYHGTIdUBlfdFYAOvbIamDQwllGxFTgNc46QGfiRIXkxJ1kLFg4x8X1KomtGI3t
VG6dMdmkMpsSMHrZn/1TZs8jFLzVZXeMSmjesQ+NwQjkW4TBg4zJ1eHvNVgM1MIp5VUnR7Yd1SmE
naiLo8RXJp6pGzG+C27CcUQhoEEBR4zhsQk2wCMFyd7pLme7MDf4aI3EMIx0ryMOB24xQ2/aCvQr
4/ySU67UMWgGcQiDxzS3ZGLBXBvlM4vMw7UY8Ggu9HDjoZwr2HvFemwKd9Pa3lOuAXj32xQ80XCO
gc96NuCJq1+6O81xuUVQJKhtn0IbJA7bZd6spJg6C5JOU+HlpFyTfUHNCkQsocpN5l507GIBwRzS
HGOccVzLPlCeFPrncH2KK4Jtbvpu3JF9EiKuYnM8QKv0gPzsp0h8gsbOrPykeo426hereJntkAQv
fSbrtsMO4Ii72ADoZi6w2BdWtSCTehrqvb6B0ZK7sGYt47GEHc+DHqhfPowmYysSYEccN3TiJ5Qc
z8IUOvGnBwJFPfVcgBwJpFf0QcFdxlN45DUfaBDpCYSBjhguM7tnQppGdjOcWlriSjriqwpE3yCG
IUdEdpd+jK+L6wtRt+8mg+zEua6/xLWKdKaN+w2TU0udIM091eYMPFt8hByMpgZOpTobc/JyGG68
QUjem7GP7jzM3RSDGRMkBI0nBhWDcJ3/FSkQZry3szHdVnapgTsLi1eY2J/STQnlyTnq9Rz0+E1u
iuD/GmHCs+5IbUNNc2x/3JpLw7+q8hU1JvVKdIgAHZvxX35YVno+AtNlnkBr3NHV/hSrhr0CoDGD
kYrCtpCNaLRjTR2O4/ITqdxpHtZAkO7UYBmLrounAbSGk7e5LbZaUt/6FflEPQJSVV+yehovDMhc
rAwH5XG331Vo1zn41a/FbDXX4FJFa2Rt97MJmLhntNlbglfQfaf605bl3ZKCjhUTjOwjZTZzrPSn
1n/9q+2MVKdDSMAg8MOIW/52ajVrQM4zIpvFMPTPfX0IoBuEWuqMWDcmgxZySMgF4D7yRwpeG7dQ
FHrPRTuMG8KRqRLgIEvBksOYYrqVQS3pt++JhaTeQhtzxfz320KlxZ6ncwRhHNClRaXE3bXTCTVE
rMKlT5bv2U3xN4prlAilZSNJDlBjR9EDUW0qUf81JZ4C3MC3VqS+M9PA4V8HPq2KjOpFIZCdfSx2
NndDLQdpwwTy/ii7mqg9MOVAuuhyTQWBexmzB41Pkx8HHQAp0GYuGvq0VgMethOYxpJb+OFvAg30
6r6JO0z9hbEYITCwpAQcXzlrA51d2KCUB/G9sRZk8yeh+UA/gFnPqdKpcW7tK+29Yu508MfOvzvY
WsDupDfxXnok9UCXrnJ8JcSXUNveD8wmFCviMWKgsHU5Qtitp3578/bf8973GHcKBUJNeYjjnWVW
Zo3uxZEqPJQvlWxCpJd5idtQy4xrfQYu0zlvyh9azZDb77iBoCj4+iqR7Qalzs8l0I6cHLpuG37o
ru3O/e4jMDVjRbCJFJkSaagyLnRUC4havSA0IIJKeHag2cZxTAf0qAx90hT3gH7RD/Wn+qEKQSqm
y0Lr2Izn1sgh2OD0SONIXTxzZzEVWOgV/IOetEcvedCPOUwGq++bsfOOY4UmEt2Idh+7kCD8lJFI
loobBhGhEBzDjAAEZVzH5jbKLZ4wVrNKXUEUAwDMb1dBj3Syhgu2iQVQjWw/nr21WS/Jm7iPNXVu
RAHMVa+8F5JRf/uHGAubY7WDEOCch56s/d++20YBfcfwGVwpzWZ6xby6crMe7XBhs4kVvZEGXke5
j5d9Mf57MB68cZM9mS8xOm+yiMGofoDIJWyNfExoJdG7iszS9SeZVzafvyN/WZk6NQlgQKE7QIXM
rp+VBjgoSgN4jY/F8Kn1LkL1YqDwk2IIvz1j6QJUyXtd8ZYbmlPeq3L7H4ypF5SG2ylN5bB4dvtV
ebqETmTwZ6cU3fBksWzXJHJP2qU0/Yp+OXtzKZwq9hz+EzHigHFQeXbGoaVxJUdy7iZEbDV2FyHs
9lgUBUB4NMNykbnp04jIsh6MaE+dGX44ZqIq+PJK5v+8Xmu+rmBFeycW9a/KoM4ea70sPABC/MZx
S4N5f3rgZmOWx9pGOyvYvwer83pKfEBxqNqGPAdzei08z2nWgT9bWCSiJZUdc8kvAsZKFrUwpp64
uS8sK2zcoFbJUfKBsugzZJUdizNU3gz0MaqBSYNicAoaXLpjkEQHtTSdTJv601epMYtUONfNxL7H
OiM89qBLHkQmU7zL+Qixtno8357mp7LILRlJEu+R1gPx+4/IAGmu8ByRsHM5O9tOzrfTL5y6g9Z/
Na/dipawK1GODPMs3qXCQPqiIDNz4t+N915T4uI60UJGgkdM+SLX32oYAVLJsqgSIhkPERKQqirK
9l7hGhCmsJ9Z06H+K4qKT56cAG5pz8sC4yLHk7DqfNM3ix5C28aYFofkXkDQc8/039ZZ9X6cMNE5
dJL2SpkfSuU33KNjZ5cld6Hxp0OttWFHgkF7V0VnOexlBuxt/oLA3wcf880Gna1bBq7zbLUtb2mQ
XaEWE5sUMYJ2e3q88pYmtlAsSpxAZ0eBWEOhCFmhIpYGbK2ITaY9cbiIR5aqdy8/oXFu4CGI+uJr
kLvWlHBYuo2IM83XawCTpbgSLu7unkP7DERrOL2rSffdlNiIyf6Vs+6IiXBgU36ECFAYTKA3w8e4
4uQBcJP5VfpQ0pX2WMTFOeCMvZxIuGQ5iRV3TCpzNaDBi5lyTNvdlay8kiTuVVvjxNiyM6eP0/tA
o6JJMzk8vAoe5ZrFZMggtTFH9O13PD29n6w9Ka+igjsyutOyb5QTu/Z6cmq4Ac3ei3DIPOeS8+7D
wBA4T5djDlbrmNE8ptejJ3/m27km8mOVBriENiSGkcu4L48EnA/SFFJ6J7Y0MBPlezZ1JssF3847
o4DTR3fBEcSPZ8q3E5bDcvd9hKS0x2CHbLSBj6heu9tUrCjv4DkUQaMyiMOvWGB1RTRTtiPoRXd/
LttGk7Nqu4Co/LxROjjcIBw5nQzBiIFFkru63v6a0ciy17v9evfwV9fmLEelwSnlycu7ldGtRWpG
RDwRYD2F+ahSxkPw0UMeK7vbFL0Iuj67lzN1CwdThcqTUat3vzBAcSGRK7zIMJJ/2LWrWTUc1/9E
ye7bFNU/CWqENoVqfG7tvi9FVYOArFnG2DcgupPf1jZdjpUtlNxyQefiBInzudbzyQIRyaPGDJnp
38+XjpTbW+ub2qyUj4Z/VJmO8KcSfzfhw3xj75V4pb2BLUUjhXn1Gig5vWszcbzXVfBlp0yq8Y3U
IJd452gxm+9LNLsLR2WVAM3ah97MWv5YakEAT2QJQesYOmB2lK7+2vu2rFr5Sgf0/mJWbRu62ct3
qizVaSUk5f4R4rRz6JQ/FkDxbEXA/8By0tIFl145qdywvhWdDnofLyaHiLbVzY+0b1+FaAzK7QvH
5EQ3ytMTaRyGfV5VcU7X7PHC7FDE1RYcFhhWsfTc2Igbr+5OHbDvsogVH3TeRO5C3JTaQulkwBV5
qJJMs3tXCcjPqebhlETAoVs7/wAEHDB/S846PgXsgoUY5x3W7l6sr7td66bDZXIs5jkl/LVTkOR/
xO+eLW1GeWca1x9MButR0M6KICApOyQrCyl9qOklsfKdz++yfBcb7qfq9hkd0POZ8/BUX6oYotGB
aguwLpo7l4wocW4Id9CMTB9+7jLavs1aZw1ucbcQCp+11ur51bFh+2VPcunJPLMm5DTZuyVoAbio
FlKWqsFmAcnic72/4DIojRnQDZcJQLxUrRhC6YP/Y8PXGwqLtHN5fGUNQlKbVQlm/80rnKVrX9cq
fNoafGiYRwCf3mJV1r/KPRQtkGy55eTLtJOYvOBRVrY2gD+O4bMincpiorYwWiepoOQaLZt32Z84
rfweA6PM1mlvwM6Igu5C++tjZluFFt7ks8e1EQyUPsrggq7OnEnrOuqIP9TlAm1M6Rap+gbvNcXF
yaERS3UUMKciMGf3V5MLrPCdTT8UbcgMYbySnyJ7bmONUg2zKDrVas3nOZhc/iLViIfxflWyYw2W
4hZcP6TR6UxKEQ2wGXWai346j/8v3mpnQh5QSKUE2KI0CypVeTA7N7hx9HU4bgkp4EB8L6YRyyjP
TVsOTOuXwo9RmE87TZ2cF0Nc3x23MaS4TIeS0s9Ty1K2YKPt5/8YqOlmNouKROrAnZepIqy1bWku
UV0HajVsmppsFtoQKsjftb51ONNuu/sfb2yltDl6EzJaaBMRpo2cAekhlBB1CjNoqUyE4aQBsntn
Ka7YrsmPHLz5DYKFyDLKYGAAWZGZEi5PRtGHgah1l7ghTLMD6n20OXlPHHnW985FGZmKe25Gk1gn
en8132N+2dP8OFztv+b+l4chEWWBNrMa/DZ3npbjkKQRJ770rn94mTOr9rofUstWMgdMR9FJ8qjq
039Lm+vzo8BtYCeezRW2dl3AMs7IRa9VioZndYjbNS6L3bDe8K8og/8bYHxTlkCAssvT5dx5uF+B
e8rq8IMLEWGfCj+iPMBSz/tMUM78JYr99VIJNXOwOMWTgyloFmag7+ZoPQyQJE8l9z73sWSvg+pe
PhZVRGvIkVs6KcnWRWaEiE9DbgZaT7/DdyjMgLZw1snf0f9ozEcOwoRuJNYvr5K2SFDktCQHww+l
czvfvBkhBSLhpVGSME5WDJPjDaXKcbiZ+LMJW/1mdlwEzz7Qs7XZp7Ev/FY9ydyYQb/bjPNA6OpO
AeSSROuwpFWlWEVH37n4rH2LLm5W/GN63bAqxbw8xPxjHkcKAQ54xXOYPfv0vNAVeIcqyJ2gNBbU
dFVtlFtB0CZ/tTn6DGapqo8ZODLav0uDlQ08cuvAaLSXuGSLDCk/bcZeQC4y/ZwXu8H0+eiUsKyY
+qzj+8cwxHZkfBM+amOsgNl/vc6ZIve8D+cIq14zeic3YYl5dT1Q18ek89vy/ktGV28lvkhniurh
tOyxzUwhU9ACfuY2VfXNjxCLFkQtkO7/UcInt7cT1WQunZvQvZwWYWgPVqgo2P4Le24scJfbCLMP
5IOn+DjL9+64Qe27Oq6neRGhHG2JY0IfH8bBIdPzG8cVKVWDRb7dG0c6BXwj8B6nDIwbUQurlSYS
/eDCqvLK+bVaUPMkAjWgNsJ31T9UYvBt3SxApVaBzZbSruR44dnHIw2x6NS/C+spb5lVGMrBp/j+
8CgT4yg8609m5B90GD8AZB7u2AjdwENGnn0aDmWuwYCxauQN2XjC7Y+sh5/ZTZcyQTlrct/Hem5H
AAD4ci6nrZGmkvsnHMmiSdCssXADxbS03vvFVndpIKGvvJZ4MT+mfwxtTwPCyIEPFlsl9zEjmKQD
WPYyhHUBXwWE5SZlIPrsIh2Sw6MUG0v9ryvJR94thVNwza3H+UhMCqOcGQFYUOgFOYrPxHiTay+r
QEHqj/B0o8rtJJ2BHQpwHNpurldc1tY7x5cxG+pg0igWSqPnVrIJQOofyVsGQbzaaNCJylu5a1lJ
TWEH/ShhkHjjhOVqh23WxJtFpgbM7ANpHt9lEb/A02lYWEltsFKS2H/FG7+TTDCiCURF+lz6piUH
/FilpejcNJh8Z1sN/TxymR/4DvluH2eftZlbzob6txG5Hp67ttUK5ZIMouojU9gasgr/deZdNAc4
+nF/+4M938AIpQHeSLnp4tHdKCZwMQLKxKlM+BbJ3/4VoEPTuTqZrbDh4p/wYtPNadG1+CR+Gtim
TKYxPOfbyjYPEQKsrYaJawZCntaGClQA/g+vmoMH2xFFljY4N4a7nng0CxuatrGwY5GcT2WXQg82
mU3/v5IDd0/p7jC9SD17mfmyjWN+7Njo/MKnF5ToZ+kZUb6UReJFleeg/M3JQ+pX3kpIOlABDrC8
hvFuqMuy1kZ8PgCkwH0fTG0w6+XF0I089vUqtSGtDBsIqewzIEbuLnu7JCenugmc2idjCRexmy0c
Z1qewK2vGityP0CobihhEybK0eOvxBMwV6OuoneChB/z8gLynEuzzBTxlN4nBisLfKv6zY4KOQn2
7mav2uuNQkX7xz8nZN27eIwmVcNi2SFZjAC1ZKVeqXAwYA0YvgaStjduU2hnCCAuAoIlFZmlQqFJ
kRlJ7u0/BaTYWcR0FenD9CHzJx93B8q2SS8cUfmIsPJrHqYNC65F4RJpI/TesQWWu1FwnPQ4CFfu
ipNjBasoTxmdgFOobO9Twv+C3Ab8hyqX9aiejyFbVD8V4/Zv6L5L1v53E9reOYoru3IBp4DUZ4gI
0wPFeHoWfucLBOWpEwEtQgGTpFlBwZ0AAuoQ+OpbvnWt9nt4/3s2eogs49wUETgDnApoS8kCEC0L
jENPej7YEwBTxBXVjkEh++GZJBVDlcaOWHt9+6IvIXT29EiApjySGjgvGYrhh3m2YdQuHDw+GIjl
1/O5mv0NXDVHLGmGaiEdCIiD0PMeQI0Bb9+ZfpF3puvmvscJ9C5WmwiqChy04Ea3htNl1Pb6Wwv+
UhIq0B9I18QFNi0LurLZsCqg0mcGNGGWyBGQAdKe/vLaak08+MSfmZrBCmO8ewc3pajo9FyZLynG
hfHiUivfuHrSvgN+27NYdPXcIvFZ4coWUfUilmyhpC0Bc9GEiR7wugEpHtTwYbELwB/VBt1SCQBG
DmGtZWk2q8xHyXfVYEvJE3uKdP2Zfd219h3hGSzYwZGta5A+4DiIPL8/ZAvxUcWryUACz3pYpr5z
T/2QrSNAvtaFbWwuA3BWmEOvIsySU9nR4H8Q7J7RJZWMr5DSKNQl6j7DnUsb+gx2bGfSoI9MmmH/
rB88YYx2yVgpupP0LYNN6JbD6lKibXCAilaNRR7zWqidGWPnCFY1fPMSeECy+ZqqG0U5ErBlAa4u
pOZWKrXRpvDUSao8q1M+DSK7GGT2fYXzRo4pscXQEToI760mWfzwBJzoPiN68d06cxakifbYzul8
AOtsHet4T4btmjsY2wz6ekXLZPp17jOJ6o9sXfYT2VRGuDBZ5Tlw66G/l0HdW0ar0U0o0ye4qHTU
bxtVSZT5GVKeaqyuj50U2X6UCmL3NWZ2yZalb2waLgifO9m4m4IlHvjtjAylApNApL4oeHMq8z9Y
SqvqWu8KszWMBzsIyibZH/knlVX7SBSTGrDt9jWJSShrqsjuiCvhEyPAxSzRB7q0LDEoa+ZNH+2t
zbrRZGVYgFzsL2bJDC2ZSctpX+feKDyRD+3+gef1WXEiwYyqfq7l9oUZhWBRHbIfLGcpcuE2lKsy
v8do9t7T0Wit/wng5HU91EmWF+cv+6Bv12VH4ljOJn2XUFyXS+Qthk4lUNmnj8VVvRXg2SzbO0W4
5MwUjgpE37sLcxTGh8p2+JzmDkYA1LtXY1+W0gqZIGw2T/yNMlteJr+UeI9+NcQ9/u9GKn/cQRVz
sWv+gkaUthdPxyXssJV1JDpWtyBb5pPsOR28ZcKdaTaMO2sQEoBrLAAY8FzHjo+FGaR3LDccePwF
3EmGDbdIv0eYmKTTnmLQtsyrOVuUwdQPdPE9kVBqaYGmzMmQoeVupJgZanAHhGCcsPFU/4YuPwT5
o62bFJYGIKJ2Wg+rzzxver2w9JPWvhc/hwusWHSYGxrMbYfux7Rwq8qI1ViNCAMeVfXKyRKdXQrV
Y11KDJWZQI0HsUeR0PoejM+KeGhhGTNCbYD0xUHTjPqDl+QkTRQ7UqBGovA2VvWuYd5ZFSc76nLK
bJUXx2cUMS72MDRwtr4myYrPeJ0AaGncCZHHH7GtK5yDhl7YDJRgKda8w75Whdbx48Ae+MiI0Qll
SpU7NvwXazFL5NyWrpo9YRiSpCXG5aQqirFY/LEbmjWtX+Q3yVAusOUt71fZVWi4+P4kUHxzELap
BNpgVMR677AEihPWBd1ie8o4E1AS6QhZGJjP+Uk+MDbiySzOV1laIC3Fdm4+R7OT4YAxGtHbA/Md
pAT/GDwNjagfkLPsypgxHI9Er7tDea478UkCh4BKHsPN3fULp9BYUmcISTDwEa2W08XSN19o+oUf
mdxBXgghFDa6N1Z/Kgm60Cam373s8v+HoBy8/uatQgPVUUHJRnR7Pt7bjoFTIJtSrhjvOHzsNzaw
DXwdmIrmsZfdRpe3eAkA3EwHotV/42LWZep+Ddbq4O2BQ8EFr0Wn0LJQGz0w6r6zMdRqP/37ZrlT
CQcChzZWgsEVi4SsGDz2rqPr8+T/CMw6fcdUnURZMJbA2z0Xcf1g2OImt1vk9G1ImS57bomn2Wbg
FalDfqWs6Wm+HuK3M7Qt/mrd+5LxcQ92bUXHcFIT1wJvJEeyIFDqwHzy3y0ctvCrpdhIta0U4vax
6vGk3eWAtBuRrXcnPnUVX/m2cZX0gqR3sHhiL8JhT+xL6BHMUM0YIOF3/S8pM/rdXo2owRYAT0Mz
taMwMVfk/FNJ6VFOhiq0z1SIzx0HE/RdDc0OVJf41vXOv3kmRwv12oHuiu/bx459hN0lkHeDlvDR
EfPcaNRejjWwGVNvb7pWs6MrqOvN+uN3HnTOtM7oKXUP9pUW7DR5dEYecJMyHgz0plmRJVXkIvkV
bc8dPM7IbfwBP3DzNqJ16LbWQYnsZv7oyIiTzecSRlnfKss1UKhgbd4AocmFTJIfck0A4OdISwmR
MdJ4LNb7PHsjDklpBQjiWw5BRam4by2CHTrRVL2n63FkA+d5TpX8AiW+X6GPOUbqBmlhJt9KNuWo
QCleXMJk/y3j2wqgzeoikLTn6ZYwd+eHaEtt3ycCyErhPcOWq+kG9CFdAJOX4Wk9uIskLDsK3ch1
ok4DKuvhm3l4JNmOJaH/CzQ9v2Qv9+2maWn0XesieNbUVNoZOr6dCi0fcnSv5CifavxLq65MqmrR
tNYK/vjM5lHPP+O59oo7xt0Xsx7GgOscpkM1zDC4UzFFhaJlks+GfikQc51IMGrTq8yep1+arsuB
Ok90KDUoK6B46mo8gybxRiIOuLKW583wIoadtgoyFsJUzk+KhkH33OAsG/1KBUm1cI3KZpbr+KkF
2chNFbsZ7XC5jGhfvARP/hiUM88xRE3/4FZV9+QEW26gxQYZerApHZ0IpUHLVAKJ+2Zmk12PVabk
FYzxwidE93LXWfu2n+zodTDDcwVGnjE8k2Yfey4RE7UrCb3MF5aqfxNLTqqmqcdGTugtcmJ7TE5w
zpzC3seTxC64ElmoODLHCrIOkyZ2IRvnb5US3t42qa53o/cA80DqAN9AFDMGW65hKubLtLwQ60N0
R+dB2DiP3WXeE23HSZQZmue3pO2FYJagjLI1bXo4XCFq5ouUnwmiuzqlD1ehg48RUe2yu6n19Iny
Fbf3BUcx6IqfZHNgKO2GDO/j49+GwLrTDEl55ZDDypThFyy4/LTDCOl8KIicd3SBysaqN77nGPia
ajFGaJrzGJwlTgeBeHepDOQtchX6qMNU7fgXCgzifwNF29rFQut4UXLjf5altac0CugedZG0PvD9
X47ovFRHDHNB3q2SuDDB1L2uULLhfNjP5+q0MzCDjSoZ2VmXu5qzOx6iTOfXatcwyVYxb65UQBEH
A4zZWLAxN0+25slxHpuT/S/eXKcFE9NgZ4rNNGEEDO7y4M/hwEM0wCW+1CYJ6Ci+qtd1J9THnsJX
3l95t7r7bamvs8sjg06jNTgCiFCk/F0dB7ow2TQxofoAKB0oT9AZbzUKl+0hsUZGIALlimJbcCXL
w38ZwUZr/yE0dpUoTqlxOT/fu5gClK2KnhAX3Eeia3rFWaqvgyyWIHZnbE5BPAzCMdYcZB/xatoN
NFeZRmcleK546eXxTkaZvkWdi/N3v+E+RbGfeQA0h9OulrHlODJQo6UPVR7ocFZ6WQ9txqm5Wu7W
4FpRLuzijtZdyg8ZFz9I+/jxyi1/VUYJulU0yD+x7Q0tkxYQQsHkihfi86kXnBeUxLUj1/JLkWMz
iaJBJD5eA427IoaRHmvqYq6xkbcjjfM1swy6sCFPP6NriKnb4zuabtdJPFLLIaxnS4DhbGZQiZAY
GKA28ERAc+1IU3aN4ORQqQK0TgU7FPiwfqKKr9HiSf8TANp7RRn0EcY8egztxQOapN7gVitBlcr4
PnAqwpRl0+iXR+PSqF9ZHoyiwEWreMIwBXjnlqf2c2wi6Cg1MtHeXKA3cnu0lft8Lkn+4p6wcIiB
Pz/4/b9J1PMm7P5eANzKO1tgUaf3Gu+5FNbi+9Gx0U77zYRMZ2uwOqSxcIK/JQDYKi21Ttjovxy+
stkktIbRE59k+9m8fN3PuLyyRzb2bUc5IffMT3VfZEEz36OXcAnEnBM+sbZePssImn9Hcf8hfb9v
29vwPS0phs8no9FVvnDxPimF/WxQG95f2PAmimh1dOMi5DqCr8rSg9LHRGPNAEfCNotxhdS/jJrf
4HtfKHT46L0jzuTnZnqGM9f09mKMd8bi1D2hyAqfNV+rsJoEIoeQRVyvt1Y+b750HEQYK9aTqGY3
dEhu9frFYulggfU/1s75I7A5Wi1Fnhdu0wnRBQm7dMzCvuoYdf9nmZj3D1KlYuMXGiR1OM4YBv1P
EUqDVRcRCUP3WIiG0Mbrbgp5N7oYc1Dn2lWXY7FrwKjWDmAyKKvCHHqZTQFeY/py/BKvg+qe+wln
+3HjaLW2QZQwGkIt6keBlzwYOX3w0LVnTkAwZnD4orW4ZObyjE0iRp5YgQ0TI6uc5G2UZX54Phh0
abBfTnNaVhzi8PbHDNEkuKOBW+sp+3pxW55ElBEy5/jpyPPFlQE3AYGJbG7vvvaSWbfcFP2CEJcp
t4z6PeFRVy9lxkGeHyBORhMVp2gTkHbzLtN1BPxpwmXMDuURkVNNLwGH/XRWdebhAfgxpDpu0CnL
MPxSVPHFpK2ENWWFFxIz/aJhKoCkddQAcdyzK+NtzjjqYeXcZ1FVb0BYstdwJteG979uKHSeY3hk
Js+mt04E3n+xzKBVjqNlLE10e2WEbWw60gsLT4mNebbuLARnigbOkfuQ8xONSMULjbk6aa78LrNi
U42zLRTux5eZO6R5WfkBMVabhIpWGVawC6lGcbJpdJidFBDXhbOfl1fYiq/yxElLJ6KPf2+0K9Wi
HOflyltKxO80wtmBMqj996jpKsp14x9SQRnwda5KbWBiC8/nbDbu6PqLuQBOvDHuq3mhfJ9IwR3V
880V6oQ17gbCe6o5NE5HQrmenJgbD2t6v8KnWOoLdaLAFQv3v6UMsWFRNIAtEI+xVst2ihjUvGB2
/rc8c+bRgnthmFjIc3Bcq4x6G2foKz7Bzt5YJblhL7Y8KZu3VLqDc6KBONZux01cS3w1Z4wtg3fg
A5VNP9EywdFkZdtsRrPAAkBU7s29UKOwXtHRdGJM6LS6ttpSx38Qh7oCOmF2FyonVDG1D/HPCgkb
mLU5RxoRvu3behCJWP/ohSdQNM4sGhcm2NGh2CvJjPU81D5cVjdTK3i/dLGl8Kk55q+c2ew0HwPH
5vpdZnjs+R+Chg3q8jglStYqH8vBOZj9J69i9VhXq6ISmB5DlFHwODBgtHXvuvxWJ7f+fnQiHn06
+9WoFfbqm+5EjwyncWatuN0EDBFZmfvZRuIPcqeCP4Ld0qcIxbfsBsR9W//DpBc1j4pQYF9CNyh9
9zSQPcWvMn701PMoh3iBzOtESAHquL/YTQwbBKlPFX/feIhzLp7J4xmfZ5pW4vu5KpWJ18g1uK/G
+PJJnHGcPWOXM8MQjUaT++i29GwNeC4TDWHbwYaJBb9z1Lsl0m6wELlgv3EjRb/3npLgexks2mr3
Avz77TsohEm4abd7Lvz/qXpzQpL5iGnoLmahRTxfuMsjWKbDmaKq97FpIl5hYNifl8JfapsvpKSY
1kq6Bbvl6v8t0dB7484EG7EWGA65Y3dc3WbGV70JkHRVJEwljIzMAHHdWqimY3eTVtwCL5bJGvJI
tkgOYL9NvznXurFnIxjQrCF//ZpWfM0UDt0W6oPGEiJWIjjpcHdprfVwRzNoJPAk7kGU2I0LzYAB
j9miwiqhHZJLM613Vxo8Ogd/FZToUFJrGQi46yRdDvXnmIfr3TgS1Gn/09hdGJMdN4giAtrTUsVs
YcIGCNl4d0+kyHaAG+pR4IpfR3eNwjKUvA7OMKLJLxh1wqgXBmLRpa1HnhLrlpMfzZ2hM68KTYqF
kE8ct2mw7tJHZK3eCbheyqCbJ/4vcb1wOonn+jUgN6H0c3Vthw5/nzjLq1WnasQI7O5PA0MUu79l
swXx+0ewDk/p0JkD/n0bX1cDdvpNqW7G4nTkei10SVF3N4TAJq5tXZShBxbmHBJzzP3h94UgYV7s
BAY4pnk8BpsaDe/Ed3bDiiJsYZcjpy34gUWxDUwTTi3//GPRm4oCgU/AI/nzXGLa4zFZlLiwDcZ9
/DvUGdoamoeLuJTtDA65npDxyoBELPLsKb4jxcI1txgDGHnx8TpEnHu8EaXFheFzxqxRaHYmXWFr
gTLqthMxWblf8eI3Nbavm+FHWb8j9aPorqWbm+qpy2XFsCNclVPwnG5dX+wEZPsmCzaFMqjphoHn
Ej5LuAPdC9o0x9bWLSoDxFc81Lk98lkom7VqvjCTPWUuAnVbFulvpghPM46yEb4+AMVnSWkOrapR
x4daoLxL94O0pl7++Ufs8QHEpMIH9kF/MFxIEphmpw50ELxi1IvK+kZLNgnVs7EI+SPh1orJSTAt
YM01UjuFvcfDj0lrWHYpjorB2ijFVmsdjY0nw0ROOx/x3afYEdVE3aCBP8NJ91KX2rAzIYTVmj8o
pXcmqDl25sH8fEErg/JFtngR72svGPFzJe+MeXATuI0xkwf+rjGLrQpMfzdijRADA/mgd/hnkdOx
JoLbWHPjbUtnJy5tu445lNQW8IddRfPIPpD6JgD7ziFHRL1HVJH0ttduJSBk/jKnSGuAiK6cg7zn
TH+BOkjPCk1rFt7BJ/YsaqZB+V0yHIIGrmFk4M9Pzersb3UGSy7J3JjTl8+aLbTcaLqzu9Usg1df
qCfHw9S94ubycdMQimlkD07ECRySlVGa+/eCeItkQcno5pbjxMt9TlOtqMYy/rjUcIeHu6SSXe5X
B6g1Z4PJjC2BmJQC2zl5PUObwASXkS3HUsFRiLjZm0kok9m4CCa25mZirvR903XDEbRlkVDxT/Fu
UrzLEqF+4HlYpm1/tjnUF+8TKBZssF6K8Ofphe7jbK9W+57HQDyVi7K5KlGx9eQ06uVnB3MWwM7F
REo2cgRXdLtbQsMidSEoUruBuXK5y5x0SjtbcQMM9SmNP1QflqmWe2Z1/O/QJL5VgKw3qBNmfrS6
wW4/Pjxlc8hgGVcEPT/o9yS7+1ko1iaCwqs9y7D79W1tsYWeajL9OP/IO7iHvIFFP7b/5DSjDvUm
L/jjAMnVysh2lEes2bBJ3DrsqBynIMTyCpVcvXZ5j/KptxwD8pfKL8FHEdSAULZD/2yN0TxuG16q
IswnKIzjVgFMX4lf4oBKe8XAuLdrzYktqUg+mnLaJHJxh4NK61rwduio6kGek+Udg6LFr/OYKXtt
15JeTJi54WCjNiV0ktZ6ikM07lE0TIkhpeg6o3e0/zByDqVWBBFvLAksq70CSBWpZ2Eov6VYsw4m
lAOVBw9IFG3aIlGy5bBDZCqSQ9rDuilrBRP5tGssvft6Tu0QeFbIwoUw3TB0XOgThs+YyFfm0vw9
h+Z50OJ7atXAXPF5C0vtm7lX/iaiiutWxtZFU/s21pONYh7kOaPkopmRiHAze0LPsQLR+E94vKXA
C4PAtSPcOSdOVkXv9Iw0SOk9Md6XJkNwVpUCnYmhLnDb3h3bU9Av7MvEAH/GxY6tQjn8k7uJyPSL
6yr037fXvpaHHMOA6F8HA9qgAZ5HOjV6c9oOUCeFYhNJSSFIiq4vW/bROPf493zaw+HR25c8IEmN
UzBqyDBcifwOVDM1/zha5jdEfJA3ivET4BPt0NR7/ibyLYAaSFPqA7gviClKmV0EGt3UgWvqWa4R
jbWsg9RHuEB+Q+QMYuuKcYTPpYue5AwDkYxTPERgbOglnBthk6/eRk6NMHKR46CGmHRFk50CGHTA
ea8BidIj+j2T/WsybbGsK3XjyrgYufhtb2IZEU4J+NfG5Nwb2o8Dn7mCA2qOovBbpxvBQlq92sbn
EFnezvTqXtYb+0/2vZU/ve+5E1QYBCgxxbCS3YyC4+LG+ww0yh0TUYVIX5PAQMN2Pue5hbyY/vQZ
rOk73Lix4QQQTYe3Ni8zD082XFA81uo/CNRxw/zJkEjmiMyYWYrViV6xRxSnf7j58qINywu/5I3m
5aiGKKwQHm2KvP1Wapni3KM7I5kXJaxVihlc1yW2o4AkDJkCLdEGTCWCw8GrVRNF5nQgCPEI6OcG
1g0Z090mqDtxXzRAn9Vqj03kHOg7djOPyqjnbk9qBQ5j4cAaH5F+kbND67bjtR2dUEoiNKf72Un8
MzPdQzyKAOiiVVLme+hd4pi9WN30n9Lk5Fo3hu3cSALqBqr/p98YD7SpOxln9NgHyYIb85j1eZfm
+vAg0rNmIH0WI8Rbx4kIlAnL4dx54csmGfyByzWPEIJQgLwsmL6t00kTsLyRv6I91KNBAXKzv4ao
sgTKlCH9iUqK3BlrJ7OP+84AfH7qaUAxi+fdJQejfnRwvQhuwpxQbYKgrRmhsHbQZSVLIBgnkKB2
uFIEogx+ydMfYBEUQhchXtg4gEnJ+6zrjdUDVniTNap9wH3+J1GNgS4k2yoKDu9xX9kSJPypLQCi
cKxdBGZ0EE39BThh+ZmYrt5tLlp2B2x9EL3wsE8yClJO/08QSP7cuKAjuIDZYGuH1b+v0/RdXeyB
4sFrLyaoWMQFLf11x+yYpcVhXKZLEfbjEPCzqoGW/nU0EWF5jk7MTaFTNSfbk5x8BJKe4YWbnvoB
RgplVt4tK0H3QJdS77QHeAMcqc5rV8HjibhZf10ZuqtYdhTjXQjvWiS9Zz6v8qBUDJU/HUnrK+1j
ciN5HX//mBKeSFBtTyR0v8u9Gf6mIsFjFdu/2cJGKxsTB2MyBSxeSBby3SxMBo/3h1N7uQYwl/5e
XtPDAGiD0FzkhluOXr3y6HysNjbNEdtoiRpLSjUelpcGhK5zb3Qp9xLP/s8hn0Q7oDdtGK+pwiMa
jrPAhAQaN1xMOvE4bPSNX5wZgLyl7jfZ0fdFSnOG+inE97zAD3iHjh9BIOkUaf0eyAIOOgFvuBUz
lhawOH8jwYE2IAlZfmWqYHx5XIEeMC+8vIhFUUPgSHDjsmYINEWwoggwLrmIuZzbptJeS0veCfln
2tTXHM4OM1Vr1ONVzYGchyUjyekbOtwDxpEl8J2tzQBw1jOaEp4QlYw6yrmhXRkOP8ptH6gsp7jU
3rQPc35omEGFw4zL5dfRTI6+yyMSHkaLMQlQqpXzTNUeN7ksYYPwhQvb57xbeI3o9iDJLEjBsX1L
i03P47vgZ2mGjZiCGZnwdExbGR3pA+EYN0hN0GvUY4nkRBrL42Rug9YSv3cJWLOYJQOP3So1usH1
qhkRqnATzLS/o71oez0K/v+R+JDuFYWiNKZWujUd3p/oJWDMd1NzjZe0RK7b4/oTTUlBHbWbQkWd
86KqNVz7F0L/ypsPU36QDFV6NbZYnNF3CXBaXghXvN8k5TSjtRGfuA57Tu5JXl7Ekmq4+Pg/J82D
wGqhShuiKsVrZZfgt8N0S1O8rchZAAuDH5N98+O+3R1vYIGrYUdkzZioNzr98p1PQvAOYZ9n3CG4
RMxsxGcop7Jtwgpm/tXTU6488t3OZKChOjyXFXNOgEkwnHgi/Hh7w3aSXea0dL0lk0wVl/QnN2C+
fHEZssWFiDxmlFsVWZvYMSKfDeV9pMZKHzQeUqKAPhMyXNdIMvMhDMMZLQD6dp169N4eVm96bay3
RFCtpfmVarqWpIZEQlvWXl4vbItLacVw5qCZPOXZFfkrqc59T7ntxXT9Kf2HJGnc3goL1MMeBAJO
czTWPzkBdthNrF3eFVp3NH+ADcqQWtzB5rpDDxDy4pG4mhvzxeYQKyyvsH0NZ1M8jXh2S+jiIx7x
aZNwrvz9M+1nwJ+thspMFDPHdJGyY1A7QMmZyY+hKPBTZoQyPt01hgCEsYc+czWFteSDmTQEclQk
jQdLTEzXdWKGZu95ptJpLcvVokjjNEzbpOeD1aWGlIXf293GLDHV43Z/uCOt9TWEiV6bG5na+AdG
nIEVFx/R5bRguSdNbdTVyZ91X/nO56CVobp3RfKs0J3gSQFC8mCd1v2u3P+VsUObQ/MP/nJ8D3Qa
THPZQwdtpoeeO0QccrdkCl5RINe64s6sKOhegeV5ldmuTSxwnmZVvdxirpzOZFcf/M9Rb8lFIlL1
+L8U5vvoPn8hzVK+6Upphn+ObsfOUZz50+5OvKcynPCy3P/AtYXc8r1K9pWveV+fATdU05osj+vT
/IWPuSGCzwwhtEkPnjLfQwFbgifdaDWgtyicEZuZf5CQo1IWeRxf2+p2TfEgg4akmydBG7mhrLUu
dJABq26Gvpsy4aL73XDBEDvW5wmgrqOMGArb/6cWpJ1drGCd4I8N7IHglJE4kRBfan/OnGx9603K
IAr/3lwaUYIuBz8G0UgKvIpbod+yEcVEl9+1Ac2M2+V2vIvS1z82tzbzRUGVsEgnbhljMDRoUZAM
FY1dfzfmgTLbrzCLMCTV//kg7ANbhJe9SboYAttUqoVIuLWe/qUeKbWU9ZsUE4ce4MMoTz3LxWtH
zRA4pCmaeYGiYDnShA4bdcqwGTeEhRpxDZfVOAiKjsIgl4jYD6Yag7e/4nZ65a+OOtxnT1LdzNb/
rK/ekW37QXUtFLR4PkvAcxtblZzLgBRbgMv1BGYSEiZ9KBhfjHsCZa0MCycxjiZLmLSyjhsCH5MK
qOZqJa3LgP2HEjZeOrCc/jm7ak8lclxoTXRFb3y1n9kf+NDw9cFu0TxQsH/aq0EOb70G0NcjHEjK
+6iknpjUb0mfoxjuok5QY0BSJgNdGswgnRCBXUR/YaoSKqmfxIPQR1nHkdPHhpaJaPg9v7JbGVgg
JxDXJTcKr/o22XJ5GgB3XxBfjQvKPuqfzP9752dKD11IsdoL6ZeBY77y72+wIhLLSokgLRWvMGvS
YijQOlZoTABtukHghbokVqhs8isszhKH9p99Ncaiq9xPN7EOhUyPUR8o3Q47XyEiNUkiknCgOrwl
OQxnll/pN+qZnzfo1Kypwe+07GQGfaif8a3a9QrF/nzFVcBu7/gQZDErETWq16pWmgqGxeM7QX2L
6sPVRBQMalYa8URGG6AzU5W/mBds2HoVg0pG90p/y+QEDO22yDwfiQ2PqoUDmrO+PGTcgEFR+5lZ
m8Xi2RpkDWJ003kTG1TO5wR9eW3xn4v28P3UK4dWed5fxkO0HIy96GygOP28VELBXVoHFIb7IiQg
1y76u/dwAgNt5fYEpeljwd0HpZIK6sS4tdpYoLoGH4eb6LPTWA6ySl124Tu0JgP/Glggtctzrt5a
jCgD6FSk8qu5/0uJTvAjpnyblEhq6Cks6YFuKIOe30Q37e6Sg7cVuMDkhQAinbK8bhh2hXZa5PdI
fGS1EpXf+d98aDq/IokUl7Q3wXZT4sA3uFILdk1oFQF2AMx7znNJ7Fc99YnvWPA1/w7Zf4vzZsry
1bTk6qbFFo6mmFluMknOIkzJP3zAHfHyvuTRCzHonsiJ/WAnpYTcdV3HwmYcSA5Uv4J0nikU4QoX
qM5E2qvi3xMNiXDmWfx7lQKXfcJW/lzTetH6R2ZNLw7S9Rckk2fpLN8sXfQl0qg5Smpn/E3HxRkR
+stnLn5uHCaWlSI5tkEUTZ6F2ao+bwigwUCcaZrsaQ5btJsqc7uxs3uFCaPUXoR+C1PzeVhCjP6d
MGaNG6DHX9rd54qfywrkqMHuHxWIQasRXXAu6LAiecxHRiYhPwqL1G17yWS0WuCFQH1Lw+vkeBiK
E/cxnsO9o/6cMqP1alcbj6qaqkmWBM9JIG1lPGG2zqiV7Y6btEw28QlwnXAKPyHpISaKlK2QR3yb
Qn8v1VsI6i5FZvfn9AbPDO+aVwpmQxxhdt5CLpTAJ9j4FqQM4AdkdXb9mreMef+7wkwWZAiK24Iu
4ViRoXqtAXzClfRmUKwHRrEZDDyi+QBCXNh3GbtIlgH/rSUKnStX7y5ml0L+NRV6xtLvCfGq7Nh9
ucQogJpPEwDahhRVr0OQ2wZL1e9o4izc5xMHY8nKtMh/Bd+MlXXHbNdjlNfAQoYD/kR/BPYqUKyA
3NRFsWUojV3EqJOao5bF9fBIwnJmllmX7S+NSUzVoD/ys4Af+K60WAyqDFkfMKf2BJH1UHyjwcbl
tbq+IRm69nR9TGyyQOJvI3gOELrHfHkv9ndGHrfkgQ+nXa6DWXc6BD+L6HgqwEH+HaExq2cRNswW
xGClDgJPBIFjHbGc+JI7mySv5WxcaSWBO225+Fux6x9uqq7QIj08GvqdinahUR/5BgGt9bSQh/aQ
XIZDEXx1JhCmWhbba/jPRxQAvZEtRaDBt9IXe2Wy2X2Hwb/qbnFSxTQ0ptxxoizZnvhfenP20pL5
lxfZwIK+rQQZ7j7G4QwA6gLKdEySDBPhDZ/kC/rZ1178wlBZjbl1+lqpBSh2GMEwlPaHF9XG0i3u
2Qwgun6mRlSJ59I6XiZTPkrDlpHroumg4zmJvTCmmESeBwUjqbVPdIZ+JHzsvwU5cVDOkPu0Vu6v
8JefN2ESINJinorJcxAezc3KnM57qtR9SPJPIveegy5EEyAcuV4wvPZcTevj1q7DXvZMNk1CMMD8
E0rENgWR0WjRu73obSGjRi9NkNKjkvwwnQGAAyZ1dYx9fjqvMjVEk/NoUvv4TzbRLPF5iaZNq+Re
GjRtZ5U+TgDeQKUJiEFBsD5HQzoCjo4UkEWJmlhL57+SYyXpklzaQ5qTzfztsWYT7JTlXCdsAg12
TekWtQljrzyOGwNR6x46R3XrOC29lWaKzfsmc3w7YEbEtjC0Pp9WXR8QjARHOIxTFyq/VhWYd5Gf
qv4plks2tsY3YSaKqiLEFW2uSksDgdpXQwpmhLRPWhVvB3CWjtSoQlqcI4U4UH81HI1k40e1TTtw
y4AcFv61igyaPdIOLrAG3ipcdoax+o7PiLUk+vm+oWuKdAyCy0yQErZYRhOzJf57uBcgLZpfohNu
dIZgdanGuaatY36I9ow4AKf6oPwndSvkeu4k0rpcPuxsIsRUb3c1JjeppUn4CSVu652hS5e2sm7i
qEEGbpalVJxNvj7ysVlbUaCKMdvC+agE/z1e3A8zvR1JIovb5iH3jgUEmxZgP3tRj7s6fdH6dFGD
ogiGNHV5TZcA2Z6Gj+1OrS7NzfyP8pxR1A6/4eLsxVsmdoj8io1Sh44ULdfATO8sOM2ocOiTvROH
GDC+YsUgA1QUua+CA3xcYnnoOTNMa08MGTD2x4COWOrI7ydSA+MjWKxCL4UlGm/LTNQlIMXm7ti1
vesbn0vCflFAhagYjJMog98UgJuwEAJl0SbS4CN/j8I/9lT/iBvgvQp48hUhiFab1nAeddOEA8En
4PZHpf+7I9uYNyDFhoGe8/lsJwWSJVidn4TnFkeNi+GomLlCy+PqKD34SSnW5sM4pgODD4Y9gMSt
GgloWreruAde0LYa/mcRw2edEkd6qH/Iskq85EmNDos2zkHGbNsluRMOE4G+Tvl4IRevPhpc+NAl
emJWjk7g12Q7vTmNwcu/hkhhjm5XaxIyuxH9tZclHh3r6HZbxgsOZX/Qf1Zdztb6iV3PldiQ05ee
9+4wqs0n9msdkzOtfhRsiQXv6ECk6TzgCejYbzCf0VXyNuRrX345y7L6cP4V+r0zoyGt7z9fLQtl
VJRelBuakytUQDs9ea9LaQ/R5U9qTqXh9+Meb7uLcXtW27qXBNxVwljAUeEK7YhfJMezRhsCxEHu
n/mQvKKjrIks3ykSVMfmhVLUN0dEM2zSbCvZMnYZiVv67L4i/EUdC53vehr6zFb8BcBtefB4XMf1
g9mtjivHG3bSJEO4ZhBSfxAlE04YciaHTlvsRDIjqkcE7l2yKvD1jNb87NZf/2rGlUQBp/Hd/P0P
3qH1jnaZoLNa4EClPswUuFCzCtcoqmO+7Wh/HYXfqcsO+b+zulqaEeI9rtr1vjIMZXICwAqqnSUX
p+1l+F5mzuC0+ggHMV0rutzbwz49cdZIh37yra/Uh2rRY/P16Rf8k5lR4dmMq8iWjZhM31CRk4xu
ubEvKOVyQSrCAHMk++MpFjMzVCm1w9LdWuoYmUKn8l6Nfbm1ewr16gkrRfLeTr9xjdKz7a0Bwn0Q
EJpZubopb/PxmVyK08yn40B/XWQ10DATYZAtQg34UywIvAhdSfHLLUT2BRAoU9YUikbRcKj3B/X7
ab4v1cZk6V21lH6/7CK5Dzal/nwDFW8L3foqMMFdGeJAyGTwum78EmsT/bvpeG5mZRe2Jn2KDlXv
SCnqq9xZn1nUE82lrjKmheHOByIhgSP/vnkdPhdg8tTJ76Gt4mGep5RqK2kE8B64altFCL+XPvgw
QQ/mIbBM2P6oXw9Z4cRBZAdt98w8YB+C11U9xcSqIND4D4qyJAYUaJUEilEXLVsdJlVyL0S8yWoJ
2/pLuUl8hFv89144CKUqL17ct2dqaao6srBjweAkCOvrBf1QzQANKgI8XN+PN/IwjlwwrGSF/zoq
2aC8HUK6Q5vtzg/VlyTZu84YjBMhrx0T5+8A7ovZTFFyofIm5a1Doa6t+i4mTdmVbGgEw85Zie4L
KBgrAIeTTlGHrQZ5lfRZ2u6crQlOf1RiK/yQ+AP+KGPSn2kmGY6RToL5+tDZ34KNCezPsOnGlksn
uVCEmjf0EasBrW88AssBaulTgS2XMipfK5+q1i9nzxTCz8EH9MeuKPR/YBBED7vDm4evP1zPRffo
68orEq5tX3P5/oiZBjUKwRyaD5o7WSkatS5qpWS2+sBLhl92Zy+r316yKYdGZiZV/c3VHB4Ug6q8
/osuZ66SLIsbGpwUDjPSzujCTBckbKWYgx2CC/jn8zWd2MnwuvH9/1trepE82oKXqpbfk4Tlhjft
TFYT7s3cEDuDdNjPiKSGCbjl+Ma3OW6K/aIenmAwOIRZChJK55RkaMQhBAm0LE3XzTTA0BtvoeIB
HVc1XvpreIVBqi9SKn274k6F1+5E8wzt7HxDKtEjZyjf5sg1rZ17L6NoKzoQfPy+gbkZS0e/HMQS
Yz0mBiQiJ3bkiSrwRKKkFpdAdsi/O6oBqsKL0SXtZMNESKfYxkqEnY+TYs4HvZLE5BCYdg3hchPz
g15pp5zCCj1sOktDnIthzzL0fvPN8xn6JRMsofl0C4dRdU9RB00AAOc4l40gxJdx1TH61pSmNxwp
aM0BAxKnNgH/6ErzcR+MklHmbjpGDhnDTeewkjDRD0aTIOXm9Zi0CBllX3vidEc1hpad2vb7vdSa
5MeboaV3QzZyclf3ox5Fz5jOtYdo4FuomKwDOUBJSaFB0ro294PXBsGpKwmMzB92mCLXCGP0Fj7c
YWyA/iYxh13fGoiwabL91AWG5ntuzjGggOhC8e3c2/spfLWm4f/QB+yxUPL//HATD/8vgns5j+W/
odVjHALvc/klJqwCcn/RWt60oNWB1GDYkxy4twvMPuXi6WVlFBYOpQ/cAY0a5eKlbblrUer43aju
9Q1I4huwAfyOHHhy4NM+UhJblpmEbdfLTOklOKP6pc9BaPUPn2wL/e+CjI2gBorUrZIucUeQ4pcF
lFerkWC6qW44goBf0VBIm72Os1MpvYPsC2O3lYf+EURNVbZ6VeHcLzBUwFYVP7wyytQT8OpuOJca
h87/dprUbsmAsBRAhaCmoTL2GlgpC/Fp8nGX9jUsGOpdpUuOKGGOjleaNvlLV6dOIhLO06D4fHHv
ILFR7ad5jjAC6V+DIMECkEfB/eKo2BkjsPfqMW5vu+m9KxtNRHVTILqsHw+1fTehxZdn427YVTq1
Sj4ifuv+ODV4ZlRNTDw7a80brLsbABwsq/eXGCvaw/r5UpJNhN1/xcfYNQ79x+wOIuMcq0WItOYX
NB2Fv5P56CkP9JXVjCmmjLT3CP0xhSAzqe9uzOi9/8Bn2/ppYQBTVNtBwxKC2t9uYkJcCFvRdj5f
56k2oOxejf5o15jRxzDP7Dcg+Cu97StbCIB8lIGA9uh5s+KdyjYZIMTBD+o7DQKppRxb8USV2134
KTijwW1FA20GjKJA2s/IdpjDdn3uHa3LruQfrB0plAtAoU99oYQF2n9sC+YbGC1p7F3o3/CV2K7U
e3yRoAWpCccTqKEdeVL7diOA8r+lne5UnHqs/Jc2q7hanA4h2f6L6TVGboRWAg7o63TEbKjkj9oF
JSoyMlixbw++ERndVuEkBh+J7Baob3wG+cBaQBguKfpraq+29TjpyR1qwmTcWr4Km9nyvhKNCENQ
k9Gmt1nSSYYhItjls6nkJFxOUjaSChuf3+FVxddjGeyuuHhK5y8dk0t6UqbPME56mIgvzq2dOB0G
y0vAlIC0GIJoHV57M9QwJg1whhQtNTF1XAIXn3wFA/6aeBD0jZR1AJ0vfj485iPb9qReLgKVX2b/
HBA59oNAKgbyLEhWTqg73Owv/9AKflK9sTvfCb9acC4Pk1RHyevjlojH5MvhpnYS9ClJd3gsxrW7
X2zgyY9fnijzssxUD9zI4vJjJ7pTR8lRJLZXWRmiEub+WeMkOFy6Y7lQ2gKOXA3dc4jrXhVg6YQO
AOxEZxaBuEbrusn09FAzl5N9FwjCmDSkhgkuP9bmugOblPvXLYTxZ8VXQOrV8D+3vANKyE2beIAM
qoT8JDWhQu00t1W66Vupq6jGoMa63B02tclhLosPUGzHFUGvEAZq3UdiW3YuZi/KtEn0FKk34Le5
Ew48dKJvjZdd97mg+tOk71yO4RfkKlSaF+JTG+pisDupJCwoESQfsiWYlbIXXdzWp04NHrtES0YG
UkUIHuk37hixrtY2x8xwvxrdfXSzrPBehgNcrgA9AOs33uzsVbF7SljSMiKskvcOQncVYc1yA83w
0VY2cimrw0iFyLJpTjW1yMkXpbPQYnHFwQedy2lE4HDc5QvDcG8DAtqY+kptAvJCQd2zCocu+0Gv
WWw3AXdbjTWgSpMALuWDCdFejBLqdx3VlvYF4BWcZtKyo1aQvVqciJkCoomSfn9CCrkNdBfhefZ2
yTdidKKUsEbju6RF8bYniSAKVdVCMoOEdMxGgV+ocPKjvnpOPre28M4Tsgt1O5WInQjGtxQl7y9q
fdkis8p2ngR0WIf9MMr1QesGzTjcqenpinL6a29T+EAAK+deKM3oXG7GzWWAiy1VsV9mgzilBepV
ykxLU/e9YzWoEldX6Ej3CZA9mBd+bS54LU/x6I2sg18b/PicHBCRgvWi4WVq4eRWmzGjC/hrMDdi
wERuC7T3tP4kmz6K14EkLqYNAJ8xBBUQ5Oik41mRpting4YJslx8hZf+qJMW2QOgmPgZAnKlY35h
4JDHxMrLJOrDHVIcXAAe7DeR37j2Ih7FdEFJQeMb/ZTL2LGJvPFqe3f6gQn3sMs10zzHFmper8uX
dDYl5JiDv9IfH0hnApIbGxksljCbHbkEh4f4E9qCS4GY1n1m8MCdfL2/tClc0Q91CEnHEElsB4Lf
NlOcfDf3bCu0QPey17/PqauAfZ0hXzJxHRHZJ7l8gFmBYNXj38JkGCVIho9JCET3wzX1MP1vYiHR
95wNBWdv4060WAIzyo0YI4EgLJYKUubMe0ZMf7yEb71jZu/aJ5mDyNfwHxd6zUMxXg4DHSccGURn
rWj8hDxQ/F85ZFKcNOJAKj3BiBjYgCzvyPIb1uptjFYaUJiQyY/WJoHox6lnKtZ6zuv5MZLEpAXs
v9vWCXHQhcOUKBc/wsubr5U7Z/2L7hgNhZjCjZaKihNt7rAYERvuO36L/l24rhuj1Lzt6rA9Gl/a
jVkERk9LEFfdlf7d69pumGBvuJMoED8S5jLpDhwajih2QfiGHiuTubdENbDt/34XsBYMm0ES6W3r
ls+YHr8KX0iWf8gXPj476GZaAR0eUhciz1tiZanfmaO9SseLU73qWoRGKBIcGM5UFcDOyeKdWqnH
6NmI1VP5EpFChawHQ5Yxw8NAhkvl2PyQp5H3R04+TuXLqBaxA3D0+OH7b37PIy+V7NtUaq7JIPtr
8lQbnSLNWO/Pq+R08h+K+8+HuKVu2eikdtjJ33CYlHYJraqCfUJS3GziF6tyRiYlJ2Zhg/TIARa9
P1pGYN6z/ioutCNsV4wXaezS1ihZ7paofdQS42bWskldfoNa3RxX9XEanFYrG0GHRxSxTLok/ybF
mL5PQldNSQ+ctTlQOxg74vplpVBuelvo8m3CJa3wBUEcIA5HQsB5wHrhRgZM7RR9U5j9NLia7wI0
isXq0dqIqLU5HZvyFYU24t6OVDp2WBcFBIrDYQ+D2WuGaE3BoMKmCQ+GUDtQKGR4wjADogjNx3fi
bEFKsJytW0USa4QyOynv1Wnvp6Le98HBoQmcuNmWHrT1zbT6q4WD/7JXt4r9OSvoX+CCCXgmikS+
1biuSbZe5nnMg11oLWM7oHWlj8Ods/INaPFOf+3zQ4WR2S1/XprYOcBjqPhOQDMW/vo9PvFoxc/J
kCjT7qmcvNK/JPzStdwCKEv2PIg5ri3o2YnVF2Eok8QPkFQTpLc7GS5zkmk5raqm9HN3Rh1Pe5RP
AUtWCCxfL4LrdyOSQaoGwRR/XW3i8J703kKmQggWjpCnvdM38bdi+J144PBvlmT2JUa2mnNO/eUg
RRvP7D10O74dhJ1YJpX9CzHJWmD4XJg5TjrTwlj72/80x1nXW46EfX5vKRt5zMb8BRJpa6gZRx57
4AD8LDgDBQPBbwjxeVc5ggsX6/s+sSOVhKCITEuzcjwNDqZ9Tu4SRbaCKov1NRm1MiCpqGLYYuUV
1pMP+cUhNDwY99c8Og98le6RK3/iyTL+H+nCVe3VVlQRtgmJr1zoCe3OEHljHAQvjENA3/fNWFcX
UmDIf8g9JG0IPBj81JKtry54tR21Udcyoox35IR8PrGAzoqPa8lsG5uXoFc5jYs4iJQ6/tj0ZjDZ
XUxG
`protect end_protected
